`timescale 1 ns / 1 ps

module wrapper_tf(

// Module IO - Clock/Reset

input wire clock,
input wire reset,

// Module IO - Bus Signals

input  wire [1:0] bus_vpf,
input  wire [3:0] bus_q,
input  wire [6:0] bus_wg,
input  wire [7:0] bus_hstr,
input  wire [3:0] bus_cpat,
input  wire [10:0] bus_ph_rpc,
input  wire [4:0] bus_th_rpc,
input  wire [5:0] bus_time,
input  wire [9:0] bus_bend,
input  wire [8:0] bus_cs,
input  wire [0:0] bus_endcap,
input  wire [2:0] bus_sector,
input  wire [0:0] bus_lat_test,
input  wire [63:0] bus_core_config,
input  wire [12:0] bus_r_in,
input  wire [0:0] bus_we,
input  wire [6:0] bus_addr,
input  wire [1:0] bus_sel,
output reg [13:0] bus_model_out,
output reg [12:0] bus_r_out,

// Module IO - Control Signals

input wire feed_in_vpf,
input wire feed_in_q,
input wire feed_in_wg,
input wire feed_in_hstr,
input wire feed_in_cpat,
input wire feed_in_ph_rpc,
input wire feed_in_th_rpc,
input wire feed_in_time,
input wire feed_in_bend,
input wire feed_in_cs,
input wire feed_in_endcap,
input wire feed_in_sector,
input wire feed_in_lat_test,
input wire feed_in_core_config,
input wire feed_in_r_in,
input wire feed_in_we,
input wire feed_in_addr,
input wire feed_in_sel,
input wire feed_out_model_out,
input wire load_out_model_out,
input wire feed_out_r_out,
input wire load_out_r_out
);


// Register/Wire Declarations

reg [1:0] reg_vpf[0:11][0:8];
reg [3:0] reg_q[0:11][0:8][0:1];
reg [6:0] reg_wg[0:5][0:8][0:1];
reg [7:0] reg_hstr[0:5][0:8][0:1];
reg [3:0] reg_cpat[0:5][0:8][0:1];
reg [10:0] reg_ph_rpc[0:5][0:8][0:1];
reg [4:0] reg_th_rpc[0:5][0:8][0:1];
reg [5:0] reg_time[0:11][0:8][0:1];
reg [9:0] reg_bend[0:11][0:8][0:1];
reg [8:0] reg_cs[0:5];
reg [0:0] reg_endcap;
reg [2:0] reg_sector;
reg [0:0] reg_lat_test;
reg [63:0] reg_core_config;
reg [12:0] reg_r_in;
reg [0:0] reg_we;
reg [6:0] reg_addr;
reg [1:0] reg_sel;
reg [13:0] reg_model_out[0:215];
reg [12:0] reg_r_out;
wire [13:0] wire_model_out[0:215];
wire [12:0] wire_r_out;

    coord_delay_tl UUT (

// IO Connections

.ap_clk(clock),
.ap_rst(reset),
.vpf_0_0_V(reg_vpf[0][0]),
.vpf_0_1_V(reg_vpf[0][1]),
.vpf_0_2_V(reg_vpf[0][2]),
.vpf_0_3_V(reg_vpf[0][3]),
.vpf_0_4_V(reg_vpf[0][4]),
.vpf_0_5_V(reg_vpf[0][5]),
.vpf_0_6_V(reg_vpf[0][6]),
.vpf_0_7_V(reg_vpf[0][7]),
.vpf_0_8_V(reg_vpf[0][8]),
.vpf_1_0_V(reg_vpf[1][0]),
.vpf_1_1_V(reg_vpf[1][1]),
.vpf_1_2_V(reg_vpf[1][2]),
.vpf_1_3_V(reg_vpf[1][3]),
.vpf_1_4_V(reg_vpf[1][4]),
.vpf_1_5_V(reg_vpf[1][5]),
.vpf_1_6_V(reg_vpf[1][6]),
.vpf_1_7_V(reg_vpf[1][7]),
.vpf_1_8_V(reg_vpf[1][8]),
.vpf_2_0_V(reg_vpf[2][0]),
.vpf_2_1_V(reg_vpf[2][1]),
.vpf_2_2_V(reg_vpf[2][2]),
.vpf_2_3_V(reg_vpf[2][3]),
.vpf_2_4_V(reg_vpf[2][4]),
.vpf_2_5_V(reg_vpf[2][5]),
.vpf_2_6_V(reg_vpf[2][6]),
.vpf_2_7_V(reg_vpf[2][7]),
.vpf_2_8_V(reg_vpf[2][8]),
.vpf_3_0_V(reg_vpf[3][0]),
.vpf_3_1_V(reg_vpf[3][1]),
.vpf_3_2_V(reg_vpf[3][2]),
.vpf_3_3_V(reg_vpf[3][3]),
.vpf_3_4_V(reg_vpf[3][4]),
.vpf_3_5_V(reg_vpf[3][5]),
.vpf_3_6_V(reg_vpf[3][6]),
.vpf_3_7_V(reg_vpf[3][7]),
.vpf_3_8_V(reg_vpf[3][8]),
.vpf_4_0_V(reg_vpf[4][0]),
.vpf_4_1_V(reg_vpf[4][1]),
.vpf_4_2_V(reg_vpf[4][2]),
.vpf_4_3_V(reg_vpf[4][3]),
.vpf_4_4_V(reg_vpf[4][4]),
.vpf_4_5_V(reg_vpf[4][5]),
.vpf_4_6_V(reg_vpf[4][6]),
.vpf_4_7_V(reg_vpf[4][7]),
.vpf_4_8_V(reg_vpf[4][8]),
.vpf_5_0_V(reg_vpf[5][0]),
.vpf_5_1_V(reg_vpf[5][1]),
.vpf_5_2_V(reg_vpf[5][2]),
.vpf_5_3_V(reg_vpf[5][3]),
.vpf_5_4_V(reg_vpf[5][4]),
.vpf_5_5_V(reg_vpf[5][5]),
.vpf_5_6_V(reg_vpf[5][6]),
.vpf_5_7_V(reg_vpf[5][7]),
.vpf_5_8_V(reg_vpf[5][8]),
.vpf_6_0_V(reg_vpf[6][0]),
.vpf_6_1_V(reg_vpf[6][1]),
.vpf_6_2_V(reg_vpf[6][2]),
.vpf_6_3_V(reg_vpf[6][3]),
.vpf_6_4_V(reg_vpf[6][4]),
.vpf_6_5_V(reg_vpf[6][5]),
.vpf_6_6_V(reg_vpf[6][6]),
.vpf_6_7_V(reg_vpf[6][7]),
.vpf_6_8_V(reg_vpf[6][8]),
.vpf_7_0_V(reg_vpf[7][0]),
.vpf_7_1_V(reg_vpf[7][1]),
.vpf_7_2_V(reg_vpf[7][2]),
.vpf_7_3_V(reg_vpf[7][3]),
.vpf_7_4_V(reg_vpf[7][4]),
.vpf_7_5_V(reg_vpf[7][5]),
.vpf_7_6_V(reg_vpf[7][6]),
.vpf_7_7_V(reg_vpf[7][7]),
.vpf_7_8_V(reg_vpf[7][8]),
.vpf_8_0_V(reg_vpf[8][0]),
.vpf_8_1_V(reg_vpf[8][1]),
.vpf_8_2_V(reg_vpf[8][2]),
.vpf_8_3_V(reg_vpf[8][3]),
.vpf_8_4_V(reg_vpf[8][4]),
.vpf_8_5_V(reg_vpf[8][5]),
.vpf_8_6_V(reg_vpf[8][6]),
.vpf_8_7_V(reg_vpf[8][7]),
.vpf_8_8_V(reg_vpf[8][8]),
.vpf_9_0_V(reg_vpf[9][0]),
.vpf_9_1_V(reg_vpf[9][1]),
.vpf_9_2_V(reg_vpf[9][2]),
.vpf_9_3_V(reg_vpf[9][3]),
.vpf_9_4_V(reg_vpf[9][4]),
.vpf_9_5_V(reg_vpf[9][5]),
.vpf_9_6_V(reg_vpf[9][6]),
.vpf_9_7_V(reg_vpf[9][7]),
.vpf_9_8_V(reg_vpf[9][8]),
.vpf_10_0_V(reg_vpf[10][0]),
.vpf_10_1_V(reg_vpf[10][1]),
.vpf_10_2_V(reg_vpf[10][2]),
.vpf_10_3_V(reg_vpf[10][3]),
.vpf_10_4_V(reg_vpf[10][4]),
.vpf_10_5_V(reg_vpf[10][5]),
.vpf_10_6_V(reg_vpf[10][6]),
.vpf_10_7_V(reg_vpf[10][7]),
.vpf_10_8_V(reg_vpf[10][8]),
.vpf_11_0_V(reg_vpf[11][0]),
.vpf_11_1_V(reg_vpf[11][1]),
.vpf_11_2_V(reg_vpf[11][2]),
.vpf_11_3_V(reg_vpf[11][3]),
.vpf_11_4_V(reg_vpf[11][4]),
.vpf_11_5_V(reg_vpf[11][5]),
.vpf_11_6_V(reg_vpf[11][6]),
.vpf_11_7_V(reg_vpf[11][7]),
.vpf_11_8_V(reg_vpf[11][8]),
.q_0_0_0_V(reg_q[0][0][0]),
.q_0_0_1_V(reg_q[0][0][1]),
.q_0_1_0_V(reg_q[0][1][0]),
.q_0_1_1_V(reg_q[0][1][1]),
.q_0_2_0_V(reg_q[0][2][0]),
.q_0_2_1_V(reg_q[0][2][1]),
.q_0_3_0_V(reg_q[0][3][0]),
.q_0_3_1_V(reg_q[0][3][1]),
.q_0_4_0_V(reg_q[0][4][0]),
.q_0_4_1_V(reg_q[0][4][1]),
.q_0_5_0_V(reg_q[0][5][0]),
.q_0_5_1_V(reg_q[0][5][1]),
.q_0_6_0_V(reg_q[0][6][0]),
.q_0_6_1_V(reg_q[0][6][1]),
.q_0_7_0_V(reg_q[0][7][0]),
.q_0_7_1_V(reg_q[0][7][1]),
.q_0_8_0_V(reg_q[0][8][0]),
.q_0_8_1_V(reg_q[0][8][1]),
.q_1_0_0_V(reg_q[1][0][0]),
.q_1_0_1_V(reg_q[1][0][1]),
.q_1_1_0_V(reg_q[1][1][0]),
.q_1_1_1_V(reg_q[1][1][1]),
.q_1_2_0_V(reg_q[1][2][0]),
.q_1_2_1_V(reg_q[1][2][1]),
.q_1_3_0_V(reg_q[1][3][0]),
.q_1_3_1_V(reg_q[1][3][1]),
.q_1_4_0_V(reg_q[1][4][0]),
.q_1_4_1_V(reg_q[1][4][1]),
.q_1_5_0_V(reg_q[1][5][0]),
.q_1_5_1_V(reg_q[1][5][1]),
.q_1_6_0_V(reg_q[1][6][0]),
.q_1_6_1_V(reg_q[1][6][1]),
.q_1_7_0_V(reg_q[1][7][0]),
.q_1_7_1_V(reg_q[1][7][1]),
.q_1_8_0_V(reg_q[1][8][0]),
.q_1_8_1_V(reg_q[1][8][1]),
.q_2_0_0_V(reg_q[2][0][0]),
.q_2_0_1_V(reg_q[2][0][1]),
.q_2_1_0_V(reg_q[2][1][0]),
.q_2_1_1_V(reg_q[2][1][1]),
.q_2_2_0_V(reg_q[2][2][0]),
.q_2_2_1_V(reg_q[2][2][1]),
.q_2_3_0_V(reg_q[2][3][0]),
.q_2_3_1_V(reg_q[2][3][1]),
.q_2_4_0_V(reg_q[2][4][0]),
.q_2_4_1_V(reg_q[2][4][1]),
.q_2_5_0_V(reg_q[2][5][0]),
.q_2_5_1_V(reg_q[2][5][1]),
.q_2_6_0_V(reg_q[2][6][0]),
.q_2_6_1_V(reg_q[2][6][1]),
.q_2_7_0_V(reg_q[2][7][0]),
.q_2_7_1_V(reg_q[2][7][1]),
.q_2_8_0_V(reg_q[2][8][0]),
.q_2_8_1_V(reg_q[2][8][1]),
.q_3_0_0_V(reg_q[3][0][0]),
.q_3_0_1_V(reg_q[3][0][1]),
.q_3_1_0_V(reg_q[3][1][0]),
.q_3_1_1_V(reg_q[3][1][1]),
.q_3_2_0_V(reg_q[3][2][0]),
.q_3_2_1_V(reg_q[3][2][1]),
.q_3_3_0_V(reg_q[3][3][0]),
.q_3_3_1_V(reg_q[3][3][1]),
.q_3_4_0_V(reg_q[3][4][0]),
.q_3_4_1_V(reg_q[3][4][1]),
.q_3_5_0_V(reg_q[3][5][0]),
.q_3_5_1_V(reg_q[3][5][1]),
.q_3_6_0_V(reg_q[3][6][0]),
.q_3_6_1_V(reg_q[3][6][1]),
.q_3_7_0_V(reg_q[3][7][0]),
.q_3_7_1_V(reg_q[3][7][1]),
.q_3_8_0_V(reg_q[3][8][0]),
.q_3_8_1_V(reg_q[3][8][1]),
.q_4_0_0_V(reg_q[4][0][0]),
.q_4_0_1_V(reg_q[4][0][1]),
.q_4_1_0_V(reg_q[4][1][0]),
.q_4_1_1_V(reg_q[4][1][1]),
.q_4_2_0_V(reg_q[4][2][0]),
.q_4_2_1_V(reg_q[4][2][1]),
.q_4_3_0_V(reg_q[4][3][0]),
.q_4_3_1_V(reg_q[4][3][1]),
.q_4_4_0_V(reg_q[4][4][0]),
.q_4_4_1_V(reg_q[4][4][1]),
.q_4_5_0_V(reg_q[4][5][0]),
.q_4_5_1_V(reg_q[4][5][1]),
.q_4_6_0_V(reg_q[4][6][0]),
.q_4_6_1_V(reg_q[4][6][1]),
.q_4_7_0_V(reg_q[4][7][0]),
.q_4_7_1_V(reg_q[4][7][1]),
.q_4_8_0_V(reg_q[4][8][0]),
.q_4_8_1_V(reg_q[4][8][1]),
.q_5_0_0_V(reg_q[5][0][0]),
.q_5_0_1_V(reg_q[5][0][1]),
.q_5_1_0_V(reg_q[5][1][0]),
.q_5_1_1_V(reg_q[5][1][1]),
.q_5_2_0_V(reg_q[5][2][0]),
.q_5_2_1_V(reg_q[5][2][1]),
.q_5_3_0_V(reg_q[5][3][0]),
.q_5_3_1_V(reg_q[5][3][1]),
.q_5_4_0_V(reg_q[5][4][0]),
.q_5_4_1_V(reg_q[5][4][1]),
.q_5_5_0_V(reg_q[5][5][0]),
.q_5_5_1_V(reg_q[5][5][1]),
.q_5_6_0_V(reg_q[5][6][0]),
.q_5_6_1_V(reg_q[5][6][1]),
.q_5_7_0_V(reg_q[5][7][0]),
.q_5_7_1_V(reg_q[5][7][1]),
.q_5_8_0_V(reg_q[5][8][0]),
.q_5_8_1_V(reg_q[5][8][1]),
.q_6_0_0_V(reg_q[6][0][0]),
.q_6_0_1_V(reg_q[6][0][1]),
.q_6_1_0_V(reg_q[6][1][0]),
.q_6_1_1_V(reg_q[6][1][1]),
.q_6_2_0_V(reg_q[6][2][0]),
.q_6_2_1_V(reg_q[6][2][1]),
.q_6_3_0_V(reg_q[6][3][0]),
.q_6_3_1_V(reg_q[6][3][1]),
.q_6_4_0_V(reg_q[6][4][0]),
.q_6_4_1_V(reg_q[6][4][1]),
.q_6_5_0_V(reg_q[6][5][0]),
.q_6_5_1_V(reg_q[6][5][1]),
.q_6_6_0_V(reg_q[6][6][0]),
.q_6_6_1_V(reg_q[6][6][1]),
.q_6_7_0_V(reg_q[6][7][0]),
.q_6_7_1_V(reg_q[6][7][1]),
.q_6_8_0_V(reg_q[6][8][0]),
.q_6_8_1_V(reg_q[6][8][1]),
.q_7_0_0_V(reg_q[7][0][0]),
.q_7_0_1_V(reg_q[7][0][1]),
.q_7_1_0_V(reg_q[7][1][0]),
.q_7_1_1_V(reg_q[7][1][1]),
.q_7_2_0_V(reg_q[7][2][0]),
.q_7_2_1_V(reg_q[7][2][1]),
.q_7_3_0_V(reg_q[7][3][0]),
.q_7_3_1_V(reg_q[7][3][1]),
.q_7_4_0_V(reg_q[7][4][0]),
.q_7_4_1_V(reg_q[7][4][1]),
.q_7_5_0_V(reg_q[7][5][0]),
.q_7_5_1_V(reg_q[7][5][1]),
.q_7_6_0_V(reg_q[7][6][0]),
.q_7_6_1_V(reg_q[7][6][1]),
.q_7_7_0_V(reg_q[7][7][0]),
.q_7_7_1_V(reg_q[7][7][1]),
.q_7_8_0_V(reg_q[7][8][0]),
.q_7_8_1_V(reg_q[7][8][1]),
.q_8_0_0_V(reg_q[8][0][0]),
.q_8_0_1_V(reg_q[8][0][1]),
.q_8_1_0_V(reg_q[8][1][0]),
.q_8_1_1_V(reg_q[8][1][1]),
.q_8_2_0_V(reg_q[8][2][0]),
.q_8_2_1_V(reg_q[8][2][1]),
.q_8_3_0_V(reg_q[8][3][0]),
.q_8_3_1_V(reg_q[8][3][1]),
.q_8_4_0_V(reg_q[8][4][0]),
.q_8_4_1_V(reg_q[8][4][1]),
.q_8_5_0_V(reg_q[8][5][0]),
.q_8_5_1_V(reg_q[8][5][1]),
.q_8_6_0_V(reg_q[8][6][0]),
.q_8_6_1_V(reg_q[8][6][1]),
.q_8_7_0_V(reg_q[8][7][0]),
.q_8_7_1_V(reg_q[8][7][1]),
.q_8_8_0_V(reg_q[8][8][0]),
.q_8_8_1_V(reg_q[8][8][1]),
.q_9_0_0_V(reg_q[9][0][0]),
.q_9_0_1_V(reg_q[9][0][1]),
.q_9_1_0_V(reg_q[9][1][0]),
.q_9_1_1_V(reg_q[9][1][1]),
.q_9_2_0_V(reg_q[9][2][0]),
.q_9_2_1_V(reg_q[9][2][1]),
.q_9_3_0_V(reg_q[9][3][0]),
.q_9_3_1_V(reg_q[9][3][1]),
.q_9_4_0_V(reg_q[9][4][0]),
.q_9_4_1_V(reg_q[9][4][1]),
.q_9_5_0_V(reg_q[9][5][0]),
.q_9_5_1_V(reg_q[9][5][1]),
.q_9_6_0_V(reg_q[9][6][0]),
.q_9_6_1_V(reg_q[9][6][1]),
.q_9_7_0_V(reg_q[9][7][0]),
.q_9_7_1_V(reg_q[9][7][1]),
.q_9_8_0_V(reg_q[9][8][0]),
.q_9_8_1_V(reg_q[9][8][1]),
.q_10_0_0_V(reg_q[10][0][0]),
.q_10_0_1_V(reg_q[10][0][1]),
.q_10_1_0_V(reg_q[10][1][0]),
.q_10_1_1_V(reg_q[10][1][1]),
.q_10_2_0_V(reg_q[10][2][0]),
.q_10_2_1_V(reg_q[10][2][1]),
.q_10_3_0_V(reg_q[10][3][0]),
.q_10_3_1_V(reg_q[10][3][1]),
.q_10_4_0_V(reg_q[10][4][0]),
.q_10_4_1_V(reg_q[10][4][1]),
.q_10_5_0_V(reg_q[10][5][0]),
.q_10_5_1_V(reg_q[10][5][1]),
.q_10_6_0_V(reg_q[10][6][0]),
.q_10_6_1_V(reg_q[10][6][1]),
.q_10_7_0_V(reg_q[10][7][0]),
.q_10_7_1_V(reg_q[10][7][1]),
.q_10_8_0_V(reg_q[10][8][0]),
.q_10_8_1_V(reg_q[10][8][1]),
.q_11_0_0_V(reg_q[11][0][0]),
.q_11_0_1_V(reg_q[11][0][1]),
.q_11_1_0_V(reg_q[11][1][0]),
.q_11_1_1_V(reg_q[11][1][1]),
.q_11_2_0_V(reg_q[11][2][0]),
.q_11_2_1_V(reg_q[11][2][1]),
.q_11_3_0_V(reg_q[11][3][0]),
.q_11_3_1_V(reg_q[11][3][1]),
.q_11_4_0_V(reg_q[11][4][0]),
.q_11_4_1_V(reg_q[11][4][1]),
.q_11_5_0_V(reg_q[11][5][0]),
.q_11_5_1_V(reg_q[11][5][1]),
.q_11_6_0_V(reg_q[11][6][0]),
.q_11_6_1_V(reg_q[11][6][1]),
.q_11_7_0_V(reg_q[11][7][0]),
.q_11_7_1_V(reg_q[11][7][1]),
.q_11_8_0_V(reg_q[11][8][0]),
.q_11_8_1_V(reg_q[11][8][1]),
.wg_0_0_0_V(reg_wg[0][0][0]),
.wg_0_0_1_V(reg_wg[0][0][1]),
.wg_0_1_0_V(reg_wg[0][1][0]),
.wg_0_1_1_V(reg_wg[0][1][1]),
.wg_0_2_0_V(reg_wg[0][2][0]),
.wg_0_2_1_V(reg_wg[0][2][1]),
.wg_0_3_0_V(reg_wg[0][3][0]),
.wg_0_3_1_V(reg_wg[0][3][1]),
.wg_0_4_0_V(reg_wg[0][4][0]),
.wg_0_4_1_V(reg_wg[0][4][1]),
.wg_0_5_0_V(reg_wg[0][5][0]),
.wg_0_5_1_V(reg_wg[0][5][1]),
.wg_0_6_0_V(reg_wg[0][6][0]),
.wg_0_6_1_V(reg_wg[0][6][1]),
.wg_0_7_0_V(reg_wg[0][7][0]),
.wg_0_7_1_V(reg_wg[0][7][1]),
.wg_0_8_0_V(reg_wg[0][8][0]),
.wg_0_8_1_V(reg_wg[0][8][1]),
.wg_1_0_0_V(reg_wg[1][0][0]),
.wg_1_0_1_V(reg_wg[1][0][1]),
.wg_1_1_0_V(reg_wg[1][1][0]),
.wg_1_1_1_V(reg_wg[1][1][1]),
.wg_1_2_0_V(reg_wg[1][2][0]),
.wg_1_2_1_V(reg_wg[1][2][1]),
.wg_1_3_0_V(reg_wg[1][3][0]),
.wg_1_3_1_V(reg_wg[1][3][1]),
.wg_1_4_0_V(reg_wg[1][4][0]),
.wg_1_4_1_V(reg_wg[1][4][1]),
.wg_1_5_0_V(reg_wg[1][5][0]),
.wg_1_5_1_V(reg_wg[1][5][1]),
.wg_1_6_0_V(reg_wg[1][6][0]),
.wg_1_6_1_V(reg_wg[1][6][1]),
.wg_1_7_0_V(reg_wg[1][7][0]),
.wg_1_7_1_V(reg_wg[1][7][1]),
.wg_1_8_0_V(reg_wg[1][8][0]),
.wg_1_8_1_V(reg_wg[1][8][1]),
.wg_2_0_0_V(reg_wg[2][0][0]),
.wg_2_0_1_V(reg_wg[2][0][1]),
.wg_2_1_0_V(reg_wg[2][1][0]),
.wg_2_1_1_V(reg_wg[2][1][1]),
.wg_2_2_0_V(reg_wg[2][2][0]),
.wg_2_2_1_V(reg_wg[2][2][1]),
.wg_2_3_0_V(reg_wg[2][3][0]),
.wg_2_3_1_V(reg_wg[2][3][1]),
.wg_2_4_0_V(reg_wg[2][4][0]),
.wg_2_4_1_V(reg_wg[2][4][1]),
.wg_2_5_0_V(reg_wg[2][5][0]),
.wg_2_5_1_V(reg_wg[2][5][1]),
.wg_2_6_0_V(reg_wg[2][6][0]),
.wg_2_6_1_V(reg_wg[2][6][1]),
.wg_2_7_0_V(reg_wg[2][7][0]),
.wg_2_7_1_V(reg_wg[2][7][1]),
.wg_2_8_0_V(reg_wg[2][8][0]),
.wg_2_8_1_V(reg_wg[2][8][1]),
.wg_3_0_0_V(reg_wg[3][0][0]),
.wg_3_0_1_V(reg_wg[3][0][1]),
.wg_3_1_0_V(reg_wg[3][1][0]),
.wg_3_1_1_V(reg_wg[3][1][1]),
.wg_3_2_0_V(reg_wg[3][2][0]),
.wg_3_2_1_V(reg_wg[3][2][1]),
.wg_3_3_0_V(reg_wg[3][3][0]),
.wg_3_3_1_V(reg_wg[3][3][1]),
.wg_3_4_0_V(reg_wg[3][4][0]),
.wg_3_4_1_V(reg_wg[3][4][1]),
.wg_3_5_0_V(reg_wg[3][5][0]),
.wg_3_5_1_V(reg_wg[3][5][1]),
.wg_3_6_0_V(reg_wg[3][6][0]),
.wg_3_6_1_V(reg_wg[3][6][1]),
.wg_3_7_0_V(reg_wg[3][7][0]),
.wg_3_7_1_V(reg_wg[3][7][1]),
.wg_3_8_0_V(reg_wg[3][8][0]),
.wg_3_8_1_V(reg_wg[3][8][1]),
.wg_4_0_0_V(reg_wg[4][0][0]),
.wg_4_0_1_V(reg_wg[4][0][1]),
.wg_4_1_0_V(reg_wg[4][1][0]),
.wg_4_1_1_V(reg_wg[4][1][1]),
.wg_4_2_0_V(reg_wg[4][2][0]),
.wg_4_2_1_V(reg_wg[4][2][1]),
.wg_4_3_0_V(reg_wg[4][3][0]),
.wg_4_3_1_V(reg_wg[4][3][1]),
.wg_4_4_0_V(reg_wg[4][4][0]),
.wg_4_4_1_V(reg_wg[4][4][1]),
.wg_4_5_0_V(reg_wg[4][5][0]),
.wg_4_5_1_V(reg_wg[4][5][1]),
.wg_4_6_0_V(reg_wg[4][6][0]),
.wg_4_6_1_V(reg_wg[4][6][1]),
.wg_4_7_0_V(reg_wg[4][7][0]),
.wg_4_7_1_V(reg_wg[4][7][1]),
.wg_4_8_0_V(reg_wg[4][8][0]),
.wg_4_8_1_V(reg_wg[4][8][1]),
.wg_5_0_0_V(reg_wg[5][0][0]),
.wg_5_0_1_V(reg_wg[5][0][1]),
.wg_5_1_0_V(reg_wg[5][1][0]),
.wg_5_1_1_V(reg_wg[5][1][1]),
.wg_5_2_0_V(reg_wg[5][2][0]),
.wg_5_2_1_V(reg_wg[5][2][1]),
.wg_5_3_0_V(reg_wg[5][3][0]),
.wg_5_3_1_V(reg_wg[5][3][1]),
.wg_5_4_0_V(reg_wg[5][4][0]),
.wg_5_4_1_V(reg_wg[5][4][1]),
.wg_5_5_0_V(reg_wg[5][5][0]),
.wg_5_5_1_V(reg_wg[5][5][1]),
.wg_5_6_0_V(reg_wg[5][6][0]),
.wg_5_6_1_V(reg_wg[5][6][1]),
.wg_5_7_0_V(reg_wg[5][7][0]),
.wg_5_7_1_V(reg_wg[5][7][1]),
.wg_5_8_0_V(reg_wg[5][8][0]),
.wg_5_8_1_V(reg_wg[5][8][1]),
.hstr_0_0_0_V(reg_hstr[0][0][0]),
.hstr_0_0_1_V(reg_hstr[0][0][1]),
.hstr_0_1_0_V(reg_hstr[0][1][0]),
.hstr_0_1_1_V(reg_hstr[0][1][1]),
.hstr_0_2_0_V(reg_hstr[0][2][0]),
.hstr_0_2_1_V(reg_hstr[0][2][1]),
.hstr_0_3_0_V(reg_hstr[0][3][0]),
.hstr_0_3_1_V(reg_hstr[0][3][1]),
.hstr_0_4_0_V(reg_hstr[0][4][0]),
.hstr_0_4_1_V(reg_hstr[0][4][1]),
.hstr_0_5_0_V(reg_hstr[0][5][0]),
.hstr_0_5_1_V(reg_hstr[0][5][1]),
.hstr_0_6_0_V(reg_hstr[0][6][0]),
.hstr_0_6_1_V(reg_hstr[0][6][1]),
.hstr_0_7_0_V(reg_hstr[0][7][0]),
.hstr_0_7_1_V(reg_hstr[0][7][1]),
.hstr_0_8_0_V(reg_hstr[0][8][0]),
.hstr_0_8_1_V(reg_hstr[0][8][1]),
.hstr_1_0_0_V(reg_hstr[1][0][0]),
.hstr_1_0_1_V(reg_hstr[1][0][1]),
.hstr_1_1_0_V(reg_hstr[1][1][0]),
.hstr_1_1_1_V(reg_hstr[1][1][1]),
.hstr_1_2_0_V(reg_hstr[1][2][0]),
.hstr_1_2_1_V(reg_hstr[1][2][1]),
.hstr_1_3_0_V(reg_hstr[1][3][0]),
.hstr_1_3_1_V(reg_hstr[1][3][1]),
.hstr_1_4_0_V(reg_hstr[1][4][0]),
.hstr_1_4_1_V(reg_hstr[1][4][1]),
.hstr_1_5_0_V(reg_hstr[1][5][0]),
.hstr_1_5_1_V(reg_hstr[1][5][1]),
.hstr_1_6_0_V(reg_hstr[1][6][0]),
.hstr_1_6_1_V(reg_hstr[1][6][1]),
.hstr_1_7_0_V(reg_hstr[1][7][0]),
.hstr_1_7_1_V(reg_hstr[1][7][1]),
.hstr_1_8_0_V(reg_hstr[1][8][0]),
.hstr_1_8_1_V(reg_hstr[1][8][1]),
.hstr_2_0_0_V(reg_hstr[2][0][0]),
.hstr_2_0_1_V(reg_hstr[2][0][1]),
.hstr_2_1_0_V(reg_hstr[2][1][0]),
.hstr_2_1_1_V(reg_hstr[2][1][1]),
.hstr_2_2_0_V(reg_hstr[2][2][0]),
.hstr_2_2_1_V(reg_hstr[2][2][1]),
.hstr_2_3_0_V(reg_hstr[2][3][0]),
.hstr_2_3_1_V(reg_hstr[2][3][1]),
.hstr_2_4_0_V(reg_hstr[2][4][0]),
.hstr_2_4_1_V(reg_hstr[2][4][1]),
.hstr_2_5_0_V(reg_hstr[2][5][0]),
.hstr_2_5_1_V(reg_hstr[2][5][1]),
.hstr_2_6_0_V(reg_hstr[2][6][0]),
.hstr_2_6_1_V(reg_hstr[2][6][1]),
.hstr_2_7_0_V(reg_hstr[2][7][0]),
.hstr_2_7_1_V(reg_hstr[2][7][1]),
.hstr_2_8_0_V(reg_hstr[2][8][0]),
.hstr_2_8_1_V(reg_hstr[2][8][1]),
.hstr_3_0_0_V(reg_hstr[3][0][0]),
.hstr_3_0_1_V(reg_hstr[3][0][1]),
.hstr_3_1_0_V(reg_hstr[3][1][0]),
.hstr_3_1_1_V(reg_hstr[3][1][1]),
.hstr_3_2_0_V(reg_hstr[3][2][0]),
.hstr_3_2_1_V(reg_hstr[3][2][1]),
.hstr_3_3_0_V(reg_hstr[3][3][0]),
.hstr_3_3_1_V(reg_hstr[3][3][1]),
.hstr_3_4_0_V(reg_hstr[3][4][0]),
.hstr_3_4_1_V(reg_hstr[3][4][1]),
.hstr_3_5_0_V(reg_hstr[3][5][0]),
.hstr_3_5_1_V(reg_hstr[3][5][1]),
.hstr_3_6_0_V(reg_hstr[3][6][0]),
.hstr_3_6_1_V(reg_hstr[3][6][1]),
.hstr_3_7_0_V(reg_hstr[3][7][0]),
.hstr_3_7_1_V(reg_hstr[3][7][1]),
.hstr_3_8_0_V(reg_hstr[3][8][0]),
.hstr_3_8_1_V(reg_hstr[3][8][1]),
.hstr_4_0_0_V(reg_hstr[4][0][0]),
.hstr_4_0_1_V(reg_hstr[4][0][1]),
.hstr_4_1_0_V(reg_hstr[4][1][0]),
.hstr_4_1_1_V(reg_hstr[4][1][1]),
.hstr_4_2_0_V(reg_hstr[4][2][0]),
.hstr_4_2_1_V(reg_hstr[4][2][1]),
.hstr_4_3_0_V(reg_hstr[4][3][0]),
.hstr_4_3_1_V(reg_hstr[4][3][1]),
.hstr_4_4_0_V(reg_hstr[4][4][0]),
.hstr_4_4_1_V(reg_hstr[4][4][1]),
.hstr_4_5_0_V(reg_hstr[4][5][0]),
.hstr_4_5_1_V(reg_hstr[4][5][1]),
.hstr_4_6_0_V(reg_hstr[4][6][0]),
.hstr_4_6_1_V(reg_hstr[4][6][1]),
.hstr_4_7_0_V(reg_hstr[4][7][0]),
.hstr_4_7_1_V(reg_hstr[4][7][1]),
.hstr_4_8_0_V(reg_hstr[4][8][0]),
.hstr_4_8_1_V(reg_hstr[4][8][1]),
.hstr_5_0_0_V(reg_hstr[5][0][0]),
.hstr_5_0_1_V(reg_hstr[5][0][1]),
.hstr_5_1_0_V(reg_hstr[5][1][0]),
.hstr_5_1_1_V(reg_hstr[5][1][1]),
.hstr_5_2_0_V(reg_hstr[5][2][0]),
.hstr_5_2_1_V(reg_hstr[5][2][1]),
.hstr_5_3_0_V(reg_hstr[5][3][0]),
.hstr_5_3_1_V(reg_hstr[5][3][1]),
.hstr_5_4_0_V(reg_hstr[5][4][0]),
.hstr_5_4_1_V(reg_hstr[5][4][1]),
.hstr_5_5_0_V(reg_hstr[5][5][0]),
.hstr_5_5_1_V(reg_hstr[5][5][1]),
.hstr_5_6_0_V(reg_hstr[5][6][0]),
.hstr_5_6_1_V(reg_hstr[5][6][1]),
.hstr_5_7_0_V(reg_hstr[5][7][0]),
.hstr_5_7_1_V(reg_hstr[5][7][1]),
.hstr_5_8_0_V(reg_hstr[5][8][0]),
.hstr_5_8_1_V(reg_hstr[5][8][1]),
.cpat_0_0_0_V(reg_cpat[0][0][0]),
.cpat_0_0_1_V(reg_cpat[0][0][1]),
.cpat_0_1_0_V(reg_cpat[0][1][0]),
.cpat_0_1_1_V(reg_cpat[0][1][1]),
.cpat_0_2_0_V(reg_cpat[0][2][0]),
.cpat_0_2_1_V(reg_cpat[0][2][1]),
.cpat_0_3_0_V(reg_cpat[0][3][0]),
.cpat_0_3_1_V(reg_cpat[0][3][1]),
.cpat_0_4_0_V(reg_cpat[0][4][0]),
.cpat_0_4_1_V(reg_cpat[0][4][1]),
.cpat_0_5_0_V(reg_cpat[0][5][0]),
.cpat_0_5_1_V(reg_cpat[0][5][1]),
.cpat_0_6_0_V(reg_cpat[0][6][0]),
.cpat_0_6_1_V(reg_cpat[0][6][1]),
.cpat_0_7_0_V(reg_cpat[0][7][0]),
.cpat_0_7_1_V(reg_cpat[0][7][1]),
.cpat_0_8_0_V(reg_cpat[0][8][0]),
.cpat_0_8_1_V(reg_cpat[0][8][1]),
.cpat_1_0_0_V(reg_cpat[1][0][0]),
.cpat_1_0_1_V(reg_cpat[1][0][1]),
.cpat_1_1_0_V(reg_cpat[1][1][0]),
.cpat_1_1_1_V(reg_cpat[1][1][1]),
.cpat_1_2_0_V(reg_cpat[1][2][0]),
.cpat_1_2_1_V(reg_cpat[1][2][1]),
.cpat_1_3_0_V(reg_cpat[1][3][0]),
.cpat_1_3_1_V(reg_cpat[1][3][1]),
.cpat_1_4_0_V(reg_cpat[1][4][0]),
.cpat_1_4_1_V(reg_cpat[1][4][1]),
.cpat_1_5_0_V(reg_cpat[1][5][0]),
.cpat_1_5_1_V(reg_cpat[1][5][1]),
.cpat_1_6_0_V(reg_cpat[1][6][0]),
.cpat_1_6_1_V(reg_cpat[1][6][1]),
.cpat_1_7_0_V(reg_cpat[1][7][0]),
.cpat_1_7_1_V(reg_cpat[1][7][1]),
.cpat_1_8_0_V(reg_cpat[1][8][0]),
.cpat_1_8_1_V(reg_cpat[1][8][1]),
.cpat_2_0_0_V(reg_cpat[2][0][0]),
.cpat_2_0_1_V(reg_cpat[2][0][1]),
.cpat_2_1_0_V(reg_cpat[2][1][0]),
.cpat_2_1_1_V(reg_cpat[2][1][1]),
.cpat_2_2_0_V(reg_cpat[2][2][0]),
.cpat_2_2_1_V(reg_cpat[2][2][1]),
.cpat_2_3_0_V(reg_cpat[2][3][0]),
.cpat_2_3_1_V(reg_cpat[2][3][1]),
.cpat_2_4_0_V(reg_cpat[2][4][0]),
.cpat_2_4_1_V(reg_cpat[2][4][1]),
.cpat_2_5_0_V(reg_cpat[2][5][0]),
.cpat_2_5_1_V(reg_cpat[2][5][1]),
.cpat_2_6_0_V(reg_cpat[2][6][0]),
.cpat_2_6_1_V(reg_cpat[2][6][1]),
.cpat_2_7_0_V(reg_cpat[2][7][0]),
.cpat_2_7_1_V(reg_cpat[2][7][1]),
.cpat_2_8_0_V(reg_cpat[2][8][0]),
.cpat_2_8_1_V(reg_cpat[2][8][1]),
.cpat_3_0_0_V(reg_cpat[3][0][0]),
.cpat_3_0_1_V(reg_cpat[3][0][1]),
.cpat_3_1_0_V(reg_cpat[3][1][0]),
.cpat_3_1_1_V(reg_cpat[3][1][1]),
.cpat_3_2_0_V(reg_cpat[3][2][0]),
.cpat_3_2_1_V(reg_cpat[3][2][1]),
.cpat_3_3_0_V(reg_cpat[3][3][0]),
.cpat_3_3_1_V(reg_cpat[3][3][1]),
.cpat_3_4_0_V(reg_cpat[3][4][0]),
.cpat_3_4_1_V(reg_cpat[3][4][1]),
.cpat_3_5_0_V(reg_cpat[3][5][0]),
.cpat_3_5_1_V(reg_cpat[3][5][1]),
.cpat_3_6_0_V(reg_cpat[3][6][0]),
.cpat_3_6_1_V(reg_cpat[3][6][1]),
.cpat_3_7_0_V(reg_cpat[3][7][0]),
.cpat_3_7_1_V(reg_cpat[3][7][1]),
.cpat_3_8_0_V(reg_cpat[3][8][0]),
.cpat_3_8_1_V(reg_cpat[3][8][1]),
.cpat_4_0_0_V(reg_cpat[4][0][0]),
.cpat_4_0_1_V(reg_cpat[4][0][1]),
.cpat_4_1_0_V(reg_cpat[4][1][0]),
.cpat_4_1_1_V(reg_cpat[4][1][1]),
.cpat_4_2_0_V(reg_cpat[4][2][0]),
.cpat_4_2_1_V(reg_cpat[4][2][1]),
.cpat_4_3_0_V(reg_cpat[4][3][0]),
.cpat_4_3_1_V(reg_cpat[4][3][1]),
.cpat_4_4_0_V(reg_cpat[4][4][0]),
.cpat_4_4_1_V(reg_cpat[4][4][1]),
.cpat_4_5_0_V(reg_cpat[4][5][0]),
.cpat_4_5_1_V(reg_cpat[4][5][1]),
.cpat_4_6_0_V(reg_cpat[4][6][0]),
.cpat_4_6_1_V(reg_cpat[4][6][1]),
.cpat_4_7_0_V(reg_cpat[4][7][0]),
.cpat_4_7_1_V(reg_cpat[4][7][1]),
.cpat_4_8_0_V(reg_cpat[4][8][0]),
.cpat_4_8_1_V(reg_cpat[4][8][1]),
.cpat_5_0_0_V(reg_cpat[5][0][0]),
.cpat_5_0_1_V(reg_cpat[5][0][1]),
.cpat_5_1_0_V(reg_cpat[5][1][0]),
.cpat_5_1_1_V(reg_cpat[5][1][1]),
.cpat_5_2_0_V(reg_cpat[5][2][0]),
.cpat_5_2_1_V(reg_cpat[5][2][1]),
.cpat_5_3_0_V(reg_cpat[5][3][0]),
.cpat_5_3_1_V(reg_cpat[5][3][1]),
.cpat_5_4_0_V(reg_cpat[5][4][0]),
.cpat_5_4_1_V(reg_cpat[5][4][1]),
.cpat_5_5_0_V(reg_cpat[5][5][0]),
.cpat_5_5_1_V(reg_cpat[5][5][1]),
.cpat_5_6_0_V(reg_cpat[5][6][0]),
.cpat_5_6_1_V(reg_cpat[5][6][1]),
.cpat_5_7_0_V(reg_cpat[5][7][0]),
.cpat_5_7_1_V(reg_cpat[5][7][1]),
.cpat_5_8_0_V(reg_cpat[5][8][0]),
.cpat_5_8_1_V(reg_cpat[5][8][1]),
.ph_rpc_0_0_0_V(reg_ph_rpc[0][0][0]),
.ph_rpc_0_0_1_V(reg_ph_rpc[0][0][1]),
.ph_rpc_0_1_0_V(reg_ph_rpc[0][1][0]),
.ph_rpc_0_1_1_V(reg_ph_rpc[0][1][1]),
.ph_rpc_0_2_0_V(reg_ph_rpc[0][2][0]),
.ph_rpc_0_2_1_V(reg_ph_rpc[0][2][1]),
.ph_rpc_0_3_0_V(reg_ph_rpc[0][3][0]),
.ph_rpc_0_3_1_V(reg_ph_rpc[0][3][1]),
.ph_rpc_0_4_0_V(reg_ph_rpc[0][4][0]),
.ph_rpc_0_4_1_V(reg_ph_rpc[0][4][1]),
.ph_rpc_0_5_0_V(reg_ph_rpc[0][5][0]),
.ph_rpc_0_5_1_V(reg_ph_rpc[0][5][1]),
.ph_rpc_0_6_0_V(reg_ph_rpc[0][6][0]),
.ph_rpc_0_6_1_V(reg_ph_rpc[0][6][1]),
.ph_rpc_0_7_0_V(reg_ph_rpc[0][7][0]),
.ph_rpc_0_7_1_V(reg_ph_rpc[0][7][1]),
.ph_rpc_0_8_0_V(reg_ph_rpc[0][8][0]),
.ph_rpc_0_8_1_V(reg_ph_rpc[0][8][1]),
.ph_rpc_1_0_0_V(reg_ph_rpc[1][0][0]),
.ph_rpc_1_0_1_V(reg_ph_rpc[1][0][1]),
.ph_rpc_1_1_0_V(reg_ph_rpc[1][1][0]),
.ph_rpc_1_1_1_V(reg_ph_rpc[1][1][1]),
.ph_rpc_1_2_0_V(reg_ph_rpc[1][2][0]),
.ph_rpc_1_2_1_V(reg_ph_rpc[1][2][1]),
.ph_rpc_1_3_0_V(reg_ph_rpc[1][3][0]),
.ph_rpc_1_3_1_V(reg_ph_rpc[1][3][1]),
.ph_rpc_1_4_0_V(reg_ph_rpc[1][4][0]),
.ph_rpc_1_4_1_V(reg_ph_rpc[1][4][1]),
.ph_rpc_1_5_0_V(reg_ph_rpc[1][5][0]),
.ph_rpc_1_5_1_V(reg_ph_rpc[1][5][1]),
.ph_rpc_1_6_0_V(reg_ph_rpc[1][6][0]),
.ph_rpc_1_6_1_V(reg_ph_rpc[1][6][1]),
.ph_rpc_1_7_0_V(reg_ph_rpc[1][7][0]),
.ph_rpc_1_7_1_V(reg_ph_rpc[1][7][1]),
.ph_rpc_1_8_0_V(reg_ph_rpc[1][8][0]),
.ph_rpc_1_8_1_V(reg_ph_rpc[1][8][1]),
.ph_rpc_2_0_0_V(reg_ph_rpc[2][0][0]),
.ph_rpc_2_0_1_V(reg_ph_rpc[2][0][1]),
.ph_rpc_2_1_0_V(reg_ph_rpc[2][1][0]),
.ph_rpc_2_1_1_V(reg_ph_rpc[2][1][1]),
.ph_rpc_2_2_0_V(reg_ph_rpc[2][2][0]),
.ph_rpc_2_2_1_V(reg_ph_rpc[2][2][1]),
.ph_rpc_2_3_0_V(reg_ph_rpc[2][3][0]),
.ph_rpc_2_3_1_V(reg_ph_rpc[2][3][1]),
.ph_rpc_2_4_0_V(reg_ph_rpc[2][4][0]),
.ph_rpc_2_4_1_V(reg_ph_rpc[2][4][1]),
.ph_rpc_2_5_0_V(reg_ph_rpc[2][5][0]),
.ph_rpc_2_5_1_V(reg_ph_rpc[2][5][1]),
.ph_rpc_2_6_0_V(reg_ph_rpc[2][6][0]),
.ph_rpc_2_6_1_V(reg_ph_rpc[2][6][1]),
.ph_rpc_2_7_0_V(reg_ph_rpc[2][7][0]),
.ph_rpc_2_7_1_V(reg_ph_rpc[2][7][1]),
.ph_rpc_2_8_0_V(reg_ph_rpc[2][8][0]),
.ph_rpc_2_8_1_V(reg_ph_rpc[2][8][1]),
.ph_rpc_3_0_0_V(reg_ph_rpc[3][0][0]),
.ph_rpc_3_0_1_V(reg_ph_rpc[3][0][1]),
.ph_rpc_3_1_0_V(reg_ph_rpc[3][1][0]),
.ph_rpc_3_1_1_V(reg_ph_rpc[3][1][1]),
.ph_rpc_3_2_0_V(reg_ph_rpc[3][2][0]),
.ph_rpc_3_2_1_V(reg_ph_rpc[3][2][1]),
.ph_rpc_3_3_0_V(reg_ph_rpc[3][3][0]),
.ph_rpc_3_3_1_V(reg_ph_rpc[3][3][1]),
.ph_rpc_3_4_0_V(reg_ph_rpc[3][4][0]),
.ph_rpc_3_4_1_V(reg_ph_rpc[3][4][1]),
.ph_rpc_3_5_0_V(reg_ph_rpc[3][5][0]),
.ph_rpc_3_5_1_V(reg_ph_rpc[3][5][1]),
.ph_rpc_3_6_0_V(reg_ph_rpc[3][6][0]),
.ph_rpc_3_6_1_V(reg_ph_rpc[3][6][1]),
.ph_rpc_3_7_0_V(reg_ph_rpc[3][7][0]),
.ph_rpc_3_7_1_V(reg_ph_rpc[3][7][1]),
.ph_rpc_3_8_0_V(reg_ph_rpc[3][8][0]),
.ph_rpc_3_8_1_V(reg_ph_rpc[3][8][1]),
.ph_rpc_4_0_0_V(reg_ph_rpc[4][0][0]),
.ph_rpc_4_0_1_V(reg_ph_rpc[4][0][1]),
.ph_rpc_4_1_0_V(reg_ph_rpc[4][1][0]),
.ph_rpc_4_1_1_V(reg_ph_rpc[4][1][1]),
.ph_rpc_4_2_0_V(reg_ph_rpc[4][2][0]),
.ph_rpc_4_2_1_V(reg_ph_rpc[4][2][1]),
.ph_rpc_4_3_0_V(reg_ph_rpc[4][3][0]),
.ph_rpc_4_3_1_V(reg_ph_rpc[4][3][1]),
.ph_rpc_4_4_0_V(reg_ph_rpc[4][4][0]),
.ph_rpc_4_4_1_V(reg_ph_rpc[4][4][1]),
.ph_rpc_4_5_0_V(reg_ph_rpc[4][5][0]),
.ph_rpc_4_5_1_V(reg_ph_rpc[4][5][1]),
.ph_rpc_4_6_0_V(reg_ph_rpc[4][6][0]),
.ph_rpc_4_6_1_V(reg_ph_rpc[4][6][1]),
.ph_rpc_4_7_0_V(reg_ph_rpc[4][7][0]),
.ph_rpc_4_7_1_V(reg_ph_rpc[4][7][1]),
.ph_rpc_4_8_0_V(reg_ph_rpc[4][8][0]),
.ph_rpc_4_8_1_V(reg_ph_rpc[4][8][1]),
.ph_rpc_5_0_0_V(reg_ph_rpc[5][0][0]),
.ph_rpc_5_0_1_V(reg_ph_rpc[5][0][1]),
.ph_rpc_5_1_0_V(reg_ph_rpc[5][1][0]),
.ph_rpc_5_1_1_V(reg_ph_rpc[5][1][1]),
.ph_rpc_5_2_0_V(reg_ph_rpc[5][2][0]),
.ph_rpc_5_2_1_V(reg_ph_rpc[5][2][1]),
.ph_rpc_5_3_0_V(reg_ph_rpc[5][3][0]),
.ph_rpc_5_3_1_V(reg_ph_rpc[5][3][1]),
.ph_rpc_5_4_0_V(reg_ph_rpc[5][4][0]),
.ph_rpc_5_4_1_V(reg_ph_rpc[5][4][1]),
.ph_rpc_5_5_0_V(reg_ph_rpc[5][5][0]),
.ph_rpc_5_5_1_V(reg_ph_rpc[5][5][1]),
.ph_rpc_5_6_0_V(reg_ph_rpc[5][6][0]),
.ph_rpc_5_6_1_V(reg_ph_rpc[5][6][1]),
.ph_rpc_5_7_0_V(reg_ph_rpc[5][7][0]),
.ph_rpc_5_7_1_V(reg_ph_rpc[5][7][1]),
.ph_rpc_5_8_0_V(reg_ph_rpc[5][8][0]),
.ph_rpc_5_8_1_V(reg_ph_rpc[5][8][1]),
.th_rpc_0_0_0_V(reg_th_rpc[0][0][0]),
.th_rpc_0_0_1_V(reg_th_rpc[0][0][1]),
.th_rpc_0_1_0_V(reg_th_rpc[0][1][0]),
.th_rpc_0_1_1_V(reg_th_rpc[0][1][1]),
.th_rpc_0_2_0_V(reg_th_rpc[0][2][0]),
.th_rpc_0_2_1_V(reg_th_rpc[0][2][1]),
.th_rpc_0_3_0_V(reg_th_rpc[0][3][0]),
.th_rpc_0_3_1_V(reg_th_rpc[0][3][1]),
.th_rpc_0_4_0_V(reg_th_rpc[0][4][0]),
.th_rpc_0_4_1_V(reg_th_rpc[0][4][1]),
.th_rpc_0_5_0_V(reg_th_rpc[0][5][0]),
.th_rpc_0_5_1_V(reg_th_rpc[0][5][1]),
.th_rpc_0_6_0_V(reg_th_rpc[0][6][0]),
.th_rpc_0_6_1_V(reg_th_rpc[0][6][1]),
.th_rpc_0_7_0_V(reg_th_rpc[0][7][0]),
.th_rpc_0_7_1_V(reg_th_rpc[0][7][1]),
.th_rpc_0_8_0_V(reg_th_rpc[0][8][0]),
.th_rpc_0_8_1_V(reg_th_rpc[0][8][1]),
.th_rpc_1_0_0_V(reg_th_rpc[1][0][0]),
.th_rpc_1_0_1_V(reg_th_rpc[1][0][1]),
.th_rpc_1_1_0_V(reg_th_rpc[1][1][0]),
.th_rpc_1_1_1_V(reg_th_rpc[1][1][1]),
.th_rpc_1_2_0_V(reg_th_rpc[1][2][0]),
.th_rpc_1_2_1_V(reg_th_rpc[1][2][1]),
.th_rpc_1_3_0_V(reg_th_rpc[1][3][0]),
.th_rpc_1_3_1_V(reg_th_rpc[1][3][1]),
.th_rpc_1_4_0_V(reg_th_rpc[1][4][0]),
.th_rpc_1_4_1_V(reg_th_rpc[1][4][1]),
.th_rpc_1_5_0_V(reg_th_rpc[1][5][0]),
.th_rpc_1_5_1_V(reg_th_rpc[1][5][1]),
.th_rpc_1_6_0_V(reg_th_rpc[1][6][0]),
.th_rpc_1_6_1_V(reg_th_rpc[1][6][1]),
.th_rpc_1_7_0_V(reg_th_rpc[1][7][0]),
.th_rpc_1_7_1_V(reg_th_rpc[1][7][1]),
.th_rpc_1_8_0_V(reg_th_rpc[1][8][0]),
.th_rpc_1_8_1_V(reg_th_rpc[1][8][1]),
.th_rpc_2_0_0_V(reg_th_rpc[2][0][0]),
.th_rpc_2_0_1_V(reg_th_rpc[2][0][1]),
.th_rpc_2_1_0_V(reg_th_rpc[2][1][0]),
.th_rpc_2_1_1_V(reg_th_rpc[2][1][1]),
.th_rpc_2_2_0_V(reg_th_rpc[2][2][0]),
.th_rpc_2_2_1_V(reg_th_rpc[2][2][1]),
.th_rpc_2_3_0_V(reg_th_rpc[2][3][0]),
.th_rpc_2_3_1_V(reg_th_rpc[2][3][1]),
.th_rpc_2_4_0_V(reg_th_rpc[2][4][0]),
.th_rpc_2_4_1_V(reg_th_rpc[2][4][1]),
.th_rpc_2_5_0_V(reg_th_rpc[2][5][0]),
.th_rpc_2_5_1_V(reg_th_rpc[2][5][1]),
.th_rpc_2_6_0_V(reg_th_rpc[2][6][0]),
.th_rpc_2_6_1_V(reg_th_rpc[2][6][1]),
.th_rpc_2_7_0_V(reg_th_rpc[2][7][0]),
.th_rpc_2_7_1_V(reg_th_rpc[2][7][1]),
.th_rpc_2_8_0_V(reg_th_rpc[2][8][0]),
.th_rpc_2_8_1_V(reg_th_rpc[2][8][1]),
.th_rpc_3_0_0_V(reg_th_rpc[3][0][0]),
.th_rpc_3_0_1_V(reg_th_rpc[3][0][1]),
.th_rpc_3_1_0_V(reg_th_rpc[3][1][0]),
.th_rpc_3_1_1_V(reg_th_rpc[3][1][1]),
.th_rpc_3_2_0_V(reg_th_rpc[3][2][0]),
.th_rpc_3_2_1_V(reg_th_rpc[3][2][1]),
.th_rpc_3_3_0_V(reg_th_rpc[3][3][0]),
.th_rpc_3_3_1_V(reg_th_rpc[3][3][1]),
.th_rpc_3_4_0_V(reg_th_rpc[3][4][0]),
.th_rpc_3_4_1_V(reg_th_rpc[3][4][1]),
.th_rpc_3_5_0_V(reg_th_rpc[3][5][0]),
.th_rpc_3_5_1_V(reg_th_rpc[3][5][1]),
.th_rpc_3_6_0_V(reg_th_rpc[3][6][0]),
.th_rpc_3_6_1_V(reg_th_rpc[3][6][1]),
.th_rpc_3_7_0_V(reg_th_rpc[3][7][0]),
.th_rpc_3_7_1_V(reg_th_rpc[3][7][1]),
.th_rpc_3_8_0_V(reg_th_rpc[3][8][0]),
.th_rpc_3_8_1_V(reg_th_rpc[3][8][1]),
.th_rpc_4_0_0_V(reg_th_rpc[4][0][0]),
.th_rpc_4_0_1_V(reg_th_rpc[4][0][1]),
.th_rpc_4_1_0_V(reg_th_rpc[4][1][0]),
.th_rpc_4_1_1_V(reg_th_rpc[4][1][1]),
.th_rpc_4_2_0_V(reg_th_rpc[4][2][0]),
.th_rpc_4_2_1_V(reg_th_rpc[4][2][1]),
.th_rpc_4_3_0_V(reg_th_rpc[4][3][0]),
.th_rpc_4_3_1_V(reg_th_rpc[4][3][1]),
.th_rpc_4_4_0_V(reg_th_rpc[4][4][0]),
.th_rpc_4_4_1_V(reg_th_rpc[4][4][1]),
.th_rpc_4_5_0_V(reg_th_rpc[4][5][0]),
.th_rpc_4_5_1_V(reg_th_rpc[4][5][1]),
.th_rpc_4_6_0_V(reg_th_rpc[4][6][0]),
.th_rpc_4_6_1_V(reg_th_rpc[4][6][1]),
.th_rpc_4_7_0_V(reg_th_rpc[4][7][0]),
.th_rpc_4_7_1_V(reg_th_rpc[4][7][1]),
.th_rpc_4_8_0_V(reg_th_rpc[4][8][0]),
.th_rpc_4_8_1_V(reg_th_rpc[4][8][1]),
.th_rpc_5_0_0_V(reg_th_rpc[5][0][0]),
.th_rpc_5_0_1_V(reg_th_rpc[5][0][1]),
.th_rpc_5_1_0_V(reg_th_rpc[5][1][0]),
.th_rpc_5_1_1_V(reg_th_rpc[5][1][1]),
.th_rpc_5_2_0_V(reg_th_rpc[5][2][0]),
.th_rpc_5_2_1_V(reg_th_rpc[5][2][1]),
.th_rpc_5_3_0_V(reg_th_rpc[5][3][0]),
.th_rpc_5_3_1_V(reg_th_rpc[5][3][1]),
.th_rpc_5_4_0_V(reg_th_rpc[5][4][0]),
.th_rpc_5_4_1_V(reg_th_rpc[5][4][1]),
.th_rpc_5_5_0_V(reg_th_rpc[5][5][0]),
.th_rpc_5_5_1_V(reg_th_rpc[5][5][1]),
.th_rpc_5_6_0_V(reg_th_rpc[5][6][0]),
.th_rpc_5_6_1_V(reg_th_rpc[5][6][1]),
.th_rpc_5_7_0_V(reg_th_rpc[5][7][0]),
.th_rpc_5_7_1_V(reg_th_rpc[5][7][1]),
.th_rpc_5_8_0_V(reg_th_rpc[5][8][0]),
.th_rpc_5_8_1_V(reg_th_rpc[5][8][1]),
.time_0_0_0_V(reg_time[0][0][0]),
.time_0_0_1_V(reg_time[0][0][1]),
.time_0_1_0_V(reg_time[0][1][0]),
.time_0_1_1_V(reg_time[0][1][1]),
.time_0_2_0_V(reg_time[0][2][0]),
.time_0_2_1_V(reg_time[0][2][1]),
.time_0_3_0_V(reg_time[0][3][0]),
.time_0_3_1_V(reg_time[0][3][1]),
.time_0_4_0_V(reg_time[0][4][0]),
.time_0_4_1_V(reg_time[0][4][1]),
.time_0_5_0_V(reg_time[0][5][0]),
.time_0_5_1_V(reg_time[0][5][1]),
.time_0_6_0_V(reg_time[0][6][0]),
.time_0_6_1_V(reg_time[0][6][1]),
.time_0_7_0_V(reg_time[0][7][0]),
.time_0_7_1_V(reg_time[0][7][1]),
.time_0_8_0_V(reg_time[0][8][0]),
.time_0_8_1_V(reg_time[0][8][1]),
.time_1_0_0_V(reg_time[1][0][0]),
.time_1_0_1_V(reg_time[1][0][1]),
.time_1_1_0_V(reg_time[1][1][0]),
.time_1_1_1_V(reg_time[1][1][1]),
.time_1_2_0_V(reg_time[1][2][0]),
.time_1_2_1_V(reg_time[1][2][1]),
.time_1_3_0_V(reg_time[1][3][0]),
.time_1_3_1_V(reg_time[1][3][1]),
.time_1_4_0_V(reg_time[1][4][0]),
.time_1_4_1_V(reg_time[1][4][1]),
.time_1_5_0_V(reg_time[1][5][0]),
.time_1_5_1_V(reg_time[1][5][1]),
.time_1_6_0_V(reg_time[1][6][0]),
.time_1_6_1_V(reg_time[1][6][1]),
.time_1_7_0_V(reg_time[1][7][0]),
.time_1_7_1_V(reg_time[1][7][1]),
.time_1_8_0_V(reg_time[1][8][0]),
.time_1_8_1_V(reg_time[1][8][1]),
.time_2_0_0_V(reg_time[2][0][0]),
.time_2_0_1_V(reg_time[2][0][1]),
.time_2_1_0_V(reg_time[2][1][0]),
.time_2_1_1_V(reg_time[2][1][1]),
.time_2_2_0_V(reg_time[2][2][0]),
.time_2_2_1_V(reg_time[2][2][1]),
.time_2_3_0_V(reg_time[2][3][0]),
.time_2_3_1_V(reg_time[2][3][1]),
.time_2_4_0_V(reg_time[2][4][0]),
.time_2_4_1_V(reg_time[2][4][1]),
.time_2_5_0_V(reg_time[2][5][0]),
.time_2_5_1_V(reg_time[2][5][1]),
.time_2_6_0_V(reg_time[2][6][0]),
.time_2_6_1_V(reg_time[2][6][1]),
.time_2_7_0_V(reg_time[2][7][0]),
.time_2_7_1_V(reg_time[2][7][1]),
.time_2_8_0_V(reg_time[2][8][0]),
.time_2_8_1_V(reg_time[2][8][1]),
.time_3_0_0_V(reg_time[3][0][0]),
.time_3_0_1_V(reg_time[3][0][1]),
.time_3_1_0_V(reg_time[3][1][0]),
.time_3_1_1_V(reg_time[3][1][1]),
.time_3_2_0_V(reg_time[3][2][0]),
.time_3_2_1_V(reg_time[3][2][1]),
.time_3_3_0_V(reg_time[3][3][0]),
.time_3_3_1_V(reg_time[3][3][1]),
.time_3_4_0_V(reg_time[3][4][0]),
.time_3_4_1_V(reg_time[3][4][1]),
.time_3_5_0_V(reg_time[3][5][0]),
.time_3_5_1_V(reg_time[3][5][1]),
.time_3_6_0_V(reg_time[3][6][0]),
.time_3_6_1_V(reg_time[3][6][1]),
.time_3_7_0_V(reg_time[3][7][0]),
.time_3_7_1_V(reg_time[3][7][1]),
.time_3_8_0_V(reg_time[3][8][0]),
.time_3_8_1_V(reg_time[3][8][1]),
.time_4_0_0_V(reg_time[4][0][0]),
.time_4_0_1_V(reg_time[4][0][1]),
.time_4_1_0_V(reg_time[4][1][0]),
.time_4_1_1_V(reg_time[4][1][1]),
.time_4_2_0_V(reg_time[4][2][0]),
.time_4_2_1_V(reg_time[4][2][1]),
.time_4_3_0_V(reg_time[4][3][0]),
.time_4_3_1_V(reg_time[4][3][1]),
.time_4_4_0_V(reg_time[4][4][0]),
.time_4_4_1_V(reg_time[4][4][1]),
.time_4_5_0_V(reg_time[4][5][0]),
.time_4_5_1_V(reg_time[4][5][1]),
.time_4_6_0_V(reg_time[4][6][0]),
.time_4_6_1_V(reg_time[4][6][1]),
.time_4_7_0_V(reg_time[4][7][0]),
.time_4_7_1_V(reg_time[4][7][1]),
.time_4_8_0_V(reg_time[4][8][0]),
.time_4_8_1_V(reg_time[4][8][1]),
.time_5_0_0_V(reg_time[5][0][0]),
.time_5_0_1_V(reg_time[5][0][1]),
.time_5_1_0_V(reg_time[5][1][0]),
.time_5_1_1_V(reg_time[5][1][1]),
.time_5_2_0_V(reg_time[5][2][0]),
.time_5_2_1_V(reg_time[5][2][1]),
.time_5_3_0_V(reg_time[5][3][0]),
.time_5_3_1_V(reg_time[5][3][1]),
.time_5_4_0_V(reg_time[5][4][0]),
.time_5_4_1_V(reg_time[5][4][1]),
.time_5_5_0_V(reg_time[5][5][0]),
.time_5_5_1_V(reg_time[5][5][1]),
.time_5_6_0_V(reg_time[5][6][0]),
.time_5_6_1_V(reg_time[5][6][1]),
.time_5_7_0_V(reg_time[5][7][0]),
.time_5_7_1_V(reg_time[5][7][1]),
.time_5_8_0_V(reg_time[5][8][0]),
.time_5_8_1_V(reg_time[5][8][1]),
.time_6_0_0_V(reg_time[6][0][0]),
.time_6_0_1_V(reg_time[6][0][1]),
.time_6_1_0_V(reg_time[6][1][0]),
.time_6_1_1_V(reg_time[6][1][1]),
.time_6_2_0_V(reg_time[6][2][0]),
.time_6_2_1_V(reg_time[6][2][1]),
.time_6_3_0_V(reg_time[6][3][0]),
.time_6_3_1_V(reg_time[6][3][1]),
.time_6_4_0_V(reg_time[6][4][0]),
.time_6_4_1_V(reg_time[6][4][1]),
.time_6_5_0_V(reg_time[6][5][0]),
.time_6_5_1_V(reg_time[6][5][1]),
.time_6_6_0_V(reg_time[6][6][0]),
.time_6_6_1_V(reg_time[6][6][1]),
.time_6_7_0_V(reg_time[6][7][0]),
.time_6_7_1_V(reg_time[6][7][1]),
.time_6_8_0_V(reg_time[6][8][0]),
.time_6_8_1_V(reg_time[6][8][1]),
.time_7_0_0_V(reg_time[7][0][0]),
.time_7_0_1_V(reg_time[7][0][1]),
.time_7_1_0_V(reg_time[7][1][0]),
.time_7_1_1_V(reg_time[7][1][1]),
.time_7_2_0_V(reg_time[7][2][0]),
.time_7_2_1_V(reg_time[7][2][1]),
.time_7_3_0_V(reg_time[7][3][0]),
.time_7_3_1_V(reg_time[7][3][1]),
.time_7_4_0_V(reg_time[7][4][0]),
.time_7_4_1_V(reg_time[7][4][1]),
.time_7_5_0_V(reg_time[7][5][0]),
.time_7_5_1_V(reg_time[7][5][1]),
.time_7_6_0_V(reg_time[7][6][0]),
.time_7_6_1_V(reg_time[7][6][1]),
.time_7_7_0_V(reg_time[7][7][0]),
.time_7_7_1_V(reg_time[7][7][1]),
.time_7_8_0_V(reg_time[7][8][0]),
.time_7_8_1_V(reg_time[7][8][1]),
.time_8_0_0_V(reg_time[8][0][0]),
.time_8_0_1_V(reg_time[8][0][1]),
.time_8_1_0_V(reg_time[8][1][0]),
.time_8_1_1_V(reg_time[8][1][1]),
.time_8_2_0_V(reg_time[8][2][0]),
.time_8_2_1_V(reg_time[8][2][1]),
.time_8_3_0_V(reg_time[8][3][0]),
.time_8_3_1_V(reg_time[8][3][1]),
.time_8_4_0_V(reg_time[8][4][0]),
.time_8_4_1_V(reg_time[8][4][1]),
.time_8_5_0_V(reg_time[8][5][0]),
.time_8_5_1_V(reg_time[8][5][1]),
.time_8_6_0_V(reg_time[8][6][0]),
.time_8_6_1_V(reg_time[8][6][1]),
.time_8_7_0_V(reg_time[8][7][0]),
.time_8_7_1_V(reg_time[8][7][1]),
.time_8_8_0_V(reg_time[8][8][0]),
.time_8_8_1_V(reg_time[8][8][1]),
.time_9_0_0_V(reg_time[9][0][0]),
.time_9_0_1_V(reg_time[9][0][1]),
.time_9_1_0_V(reg_time[9][1][0]),
.time_9_1_1_V(reg_time[9][1][1]),
.time_9_2_0_V(reg_time[9][2][0]),
.time_9_2_1_V(reg_time[9][2][1]),
.time_9_3_0_V(reg_time[9][3][0]),
.time_9_3_1_V(reg_time[9][3][1]),
.time_9_4_0_V(reg_time[9][4][0]),
.time_9_4_1_V(reg_time[9][4][1]),
.time_9_5_0_V(reg_time[9][5][0]),
.time_9_5_1_V(reg_time[9][5][1]),
.time_9_6_0_V(reg_time[9][6][0]),
.time_9_6_1_V(reg_time[9][6][1]),
.time_9_7_0_V(reg_time[9][7][0]),
.time_9_7_1_V(reg_time[9][7][1]),
.time_9_8_0_V(reg_time[9][8][0]),
.time_9_8_1_V(reg_time[9][8][1]),
.time_10_0_0_V(reg_time[10][0][0]),
.time_10_0_1_V(reg_time[10][0][1]),
.time_10_1_0_V(reg_time[10][1][0]),
.time_10_1_1_V(reg_time[10][1][1]),
.time_10_2_0_V(reg_time[10][2][0]),
.time_10_2_1_V(reg_time[10][2][1]),
.time_10_3_0_V(reg_time[10][3][0]),
.time_10_3_1_V(reg_time[10][3][1]),
.time_10_4_0_V(reg_time[10][4][0]),
.time_10_4_1_V(reg_time[10][4][1]),
.time_10_5_0_V(reg_time[10][5][0]),
.time_10_5_1_V(reg_time[10][5][1]),
.time_10_6_0_V(reg_time[10][6][0]),
.time_10_6_1_V(reg_time[10][6][1]),
.time_10_7_0_V(reg_time[10][7][0]),
.time_10_7_1_V(reg_time[10][7][1]),
.time_10_8_0_V(reg_time[10][8][0]),
.time_10_8_1_V(reg_time[10][8][1]),
.time_11_0_0_V(reg_time[11][0][0]),
.time_11_0_1_V(reg_time[11][0][1]),
.time_11_1_0_V(reg_time[11][1][0]),
.time_11_1_1_V(reg_time[11][1][1]),
.time_11_2_0_V(reg_time[11][2][0]),
.time_11_2_1_V(reg_time[11][2][1]),
.time_11_3_0_V(reg_time[11][3][0]),
.time_11_3_1_V(reg_time[11][3][1]),
.time_11_4_0_V(reg_time[11][4][0]),
.time_11_4_1_V(reg_time[11][4][1]),
.time_11_5_0_V(reg_time[11][5][0]),
.time_11_5_1_V(reg_time[11][5][1]),
.time_11_6_0_V(reg_time[11][6][0]),
.time_11_6_1_V(reg_time[11][6][1]),
.time_11_7_0_V(reg_time[11][7][0]),
.time_11_7_1_V(reg_time[11][7][1]),
.time_11_8_0_V(reg_time[11][8][0]),
.time_11_8_1_V(reg_time[11][8][1]),
.bend_0_0_0_V(reg_bend[0][0][0]),
.bend_0_0_1_V(reg_bend[0][0][1]),
.bend_0_1_0_V(reg_bend[0][1][0]),
.bend_0_1_1_V(reg_bend[0][1][1]),
.bend_0_2_0_V(reg_bend[0][2][0]),
.bend_0_2_1_V(reg_bend[0][2][1]),
.bend_0_3_0_V(reg_bend[0][3][0]),
.bend_0_3_1_V(reg_bend[0][3][1]),
.bend_0_4_0_V(reg_bend[0][4][0]),
.bend_0_4_1_V(reg_bend[0][4][1]),
.bend_0_5_0_V(reg_bend[0][5][0]),
.bend_0_5_1_V(reg_bend[0][5][1]),
.bend_0_6_0_V(reg_bend[0][6][0]),
.bend_0_6_1_V(reg_bend[0][6][1]),
.bend_0_7_0_V(reg_bend[0][7][0]),
.bend_0_7_1_V(reg_bend[0][7][1]),
.bend_0_8_0_V(reg_bend[0][8][0]),
.bend_0_8_1_V(reg_bend[0][8][1]),
.bend_1_0_0_V(reg_bend[1][0][0]),
.bend_1_0_1_V(reg_bend[1][0][1]),
.bend_1_1_0_V(reg_bend[1][1][0]),
.bend_1_1_1_V(reg_bend[1][1][1]),
.bend_1_2_0_V(reg_bend[1][2][0]),
.bend_1_2_1_V(reg_bend[1][2][1]),
.bend_1_3_0_V(reg_bend[1][3][0]),
.bend_1_3_1_V(reg_bend[1][3][1]),
.bend_1_4_0_V(reg_bend[1][4][0]),
.bend_1_4_1_V(reg_bend[1][4][1]),
.bend_1_5_0_V(reg_bend[1][5][0]),
.bend_1_5_1_V(reg_bend[1][5][1]),
.bend_1_6_0_V(reg_bend[1][6][0]),
.bend_1_6_1_V(reg_bend[1][6][1]),
.bend_1_7_0_V(reg_bend[1][7][0]),
.bend_1_7_1_V(reg_bend[1][7][1]),
.bend_1_8_0_V(reg_bend[1][8][0]),
.bend_1_8_1_V(reg_bend[1][8][1]),
.bend_2_0_0_V(reg_bend[2][0][0]),
.bend_2_0_1_V(reg_bend[2][0][1]),
.bend_2_1_0_V(reg_bend[2][1][0]),
.bend_2_1_1_V(reg_bend[2][1][1]),
.bend_2_2_0_V(reg_bend[2][2][0]),
.bend_2_2_1_V(reg_bend[2][2][1]),
.bend_2_3_0_V(reg_bend[2][3][0]),
.bend_2_3_1_V(reg_bend[2][3][1]),
.bend_2_4_0_V(reg_bend[2][4][0]),
.bend_2_4_1_V(reg_bend[2][4][1]),
.bend_2_5_0_V(reg_bend[2][5][0]),
.bend_2_5_1_V(reg_bend[2][5][1]),
.bend_2_6_0_V(reg_bend[2][6][0]),
.bend_2_6_1_V(reg_bend[2][6][1]),
.bend_2_7_0_V(reg_bend[2][7][0]),
.bend_2_7_1_V(reg_bend[2][7][1]),
.bend_2_8_0_V(reg_bend[2][8][0]),
.bend_2_8_1_V(reg_bend[2][8][1]),
.bend_3_0_0_V(reg_bend[3][0][0]),
.bend_3_0_1_V(reg_bend[3][0][1]),
.bend_3_1_0_V(reg_bend[3][1][0]),
.bend_3_1_1_V(reg_bend[3][1][1]),
.bend_3_2_0_V(reg_bend[3][2][0]),
.bend_3_2_1_V(reg_bend[3][2][1]),
.bend_3_3_0_V(reg_bend[3][3][0]),
.bend_3_3_1_V(reg_bend[3][3][1]),
.bend_3_4_0_V(reg_bend[3][4][0]),
.bend_3_4_1_V(reg_bend[3][4][1]),
.bend_3_5_0_V(reg_bend[3][5][0]),
.bend_3_5_1_V(reg_bend[3][5][1]),
.bend_3_6_0_V(reg_bend[3][6][0]),
.bend_3_6_1_V(reg_bend[3][6][1]),
.bend_3_7_0_V(reg_bend[3][7][0]),
.bend_3_7_1_V(reg_bend[3][7][1]),
.bend_3_8_0_V(reg_bend[3][8][0]),
.bend_3_8_1_V(reg_bend[3][8][1]),
.bend_4_0_0_V(reg_bend[4][0][0]),
.bend_4_0_1_V(reg_bend[4][0][1]),
.bend_4_1_0_V(reg_bend[4][1][0]),
.bend_4_1_1_V(reg_bend[4][1][1]),
.bend_4_2_0_V(reg_bend[4][2][0]),
.bend_4_2_1_V(reg_bend[4][2][1]),
.bend_4_3_0_V(reg_bend[4][3][0]),
.bend_4_3_1_V(reg_bend[4][3][1]),
.bend_4_4_0_V(reg_bend[4][4][0]),
.bend_4_4_1_V(reg_bend[4][4][1]),
.bend_4_5_0_V(reg_bend[4][5][0]),
.bend_4_5_1_V(reg_bend[4][5][1]),
.bend_4_6_0_V(reg_bend[4][6][0]),
.bend_4_6_1_V(reg_bend[4][6][1]),
.bend_4_7_0_V(reg_bend[4][7][0]),
.bend_4_7_1_V(reg_bend[4][7][1]),
.bend_4_8_0_V(reg_bend[4][8][0]),
.bend_4_8_1_V(reg_bend[4][8][1]),
.bend_5_0_0_V(reg_bend[5][0][0]),
.bend_5_0_1_V(reg_bend[5][0][1]),
.bend_5_1_0_V(reg_bend[5][1][0]),
.bend_5_1_1_V(reg_bend[5][1][1]),
.bend_5_2_0_V(reg_bend[5][2][0]),
.bend_5_2_1_V(reg_bend[5][2][1]),
.bend_5_3_0_V(reg_bend[5][3][0]),
.bend_5_3_1_V(reg_bend[5][3][1]),
.bend_5_4_0_V(reg_bend[5][4][0]),
.bend_5_4_1_V(reg_bend[5][4][1]),
.bend_5_5_0_V(reg_bend[5][5][0]),
.bend_5_5_1_V(reg_bend[5][5][1]),
.bend_5_6_0_V(reg_bend[5][6][0]),
.bend_5_6_1_V(reg_bend[5][6][1]),
.bend_5_7_0_V(reg_bend[5][7][0]),
.bend_5_7_1_V(reg_bend[5][7][1]),
.bend_5_8_0_V(reg_bend[5][8][0]),
.bend_5_8_1_V(reg_bend[5][8][1]),
.bend_6_0_0_V(reg_bend[6][0][0]),
.bend_6_0_1_V(reg_bend[6][0][1]),
.bend_6_1_0_V(reg_bend[6][1][0]),
.bend_6_1_1_V(reg_bend[6][1][1]),
.bend_6_2_0_V(reg_bend[6][2][0]),
.bend_6_2_1_V(reg_bend[6][2][1]),
.bend_6_3_0_V(reg_bend[6][3][0]),
.bend_6_3_1_V(reg_bend[6][3][1]),
.bend_6_4_0_V(reg_bend[6][4][0]),
.bend_6_4_1_V(reg_bend[6][4][1]),
.bend_6_5_0_V(reg_bend[6][5][0]),
.bend_6_5_1_V(reg_bend[6][5][1]),
.bend_6_6_0_V(reg_bend[6][6][0]),
.bend_6_6_1_V(reg_bend[6][6][1]),
.bend_6_7_0_V(reg_bend[6][7][0]),
.bend_6_7_1_V(reg_bend[6][7][1]),
.bend_6_8_0_V(reg_bend[6][8][0]),
.bend_6_8_1_V(reg_bend[6][8][1]),
.bend_7_0_0_V(reg_bend[7][0][0]),
.bend_7_0_1_V(reg_bend[7][0][1]),
.bend_7_1_0_V(reg_bend[7][1][0]),
.bend_7_1_1_V(reg_bend[7][1][1]),
.bend_7_2_0_V(reg_bend[7][2][0]),
.bend_7_2_1_V(reg_bend[7][2][1]),
.bend_7_3_0_V(reg_bend[7][3][0]),
.bend_7_3_1_V(reg_bend[7][3][1]),
.bend_7_4_0_V(reg_bend[7][4][0]),
.bend_7_4_1_V(reg_bend[7][4][1]),
.bend_7_5_0_V(reg_bend[7][5][0]),
.bend_7_5_1_V(reg_bend[7][5][1]),
.bend_7_6_0_V(reg_bend[7][6][0]),
.bend_7_6_1_V(reg_bend[7][6][1]),
.bend_7_7_0_V(reg_bend[7][7][0]),
.bend_7_7_1_V(reg_bend[7][7][1]),
.bend_7_8_0_V(reg_bend[7][8][0]),
.bend_7_8_1_V(reg_bend[7][8][1]),
.bend_8_0_0_V(reg_bend[8][0][0]),
.bend_8_0_1_V(reg_bend[8][0][1]),
.bend_8_1_0_V(reg_bend[8][1][0]),
.bend_8_1_1_V(reg_bend[8][1][1]),
.bend_8_2_0_V(reg_bend[8][2][0]),
.bend_8_2_1_V(reg_bend[8][2][1]),
.bend_8_3_0_V(reg_bend[8][3][0]),
.bend_8_3_1_V(reg_bend[8][3][1]),
.bend_8_4_0_V(reg_bend[8][4][0]),
.bend_8_4_1_V(reg_bend[8][4][1]),
.bend_8_5_0_V(reg_bend[8][5][0]),
.bend_8_5_1_V(reg_bend[8][5][1]),
.bend_8_6_0_V(reg_bend[8][6][0]),
.bend_8_6_1_V(reg_bend[8][6][1]),
.bend_8_7_0_V(reg_bend[8][7][0]),
.bend_8_7_1_V(reg_bend[8][7][1]),
.bend_8_8_0_V(reg_bend[8][8][0]),
.bend_8_8_1_V(reg_bend[8][8][1]),
.bend_9_0_0_V(reg_bend[9][0][0]),
.bend_9_0_1_V(reg_bend[9][0][1]),
.bend_9_1_0_V(reg_bend[9][1][0]),
.bend_9_1_1_V(reg_bend[9][1][1]),
.bend_9_2_0_V(reg_bend[9][2][0]),
.bend_9_2_1_V(reg_bend[9][2][1]),
.bend_9_3_0_V(reg_bend[9][3][0]),
.bend_9_3_1_V(reg_bend[9][3][1]),
.bend_9_4_0_V(reg_bend[9][4][0]),
.bend_9_4_1_V(reg_bend[9][4][1]),
.bend_9_5_0_V(reg_bend[9][5][0]),
.bend_9_5_1_V(reg_bend[9][5][1]),
.bend_9_6_0_V(reg_bend[9][6][0]),
.bend_9_6_1_V(reg_bend[9][6][1]),
.bend_9_7_0_V(reg_bend[9][7][0]),
.bend_9_7_1_V(reg_bend[9][7][1]),
.bend_9_8_0_V(reg_bend[9][8][0]),
.bend_9_8_1_V(reg_bend[9][8][1]),
.bend_10_0_0_V(reg_bend[10][0][0]),
.bend_10_0_1_V(reg_bend[10][0][1]),
.bend_10_1_0_V(reg_bend[10][1][0]),
.bend_10_1_1_V(reg_bend[10][1][1]),
.bend_10_2_0_V(reg_bend[10][2][0]),
.bend_10_2_1_V(reg_bend[10][2][1]),
.bend_10_3_0_V(reg_bend[10][3][0]),
.bend_10_3_1_V(reg_bend[10][3][1]),
.bend_10_4_0_V(reg_bend[10][4][0]),
.bend_10_4_1_V(reg_bend[10][4][1]),
.bend_10_5_0_V(reg_bend[10][5][0]),
.bend_10_5_1_V(reg_bend[10][5][1]),
.bend_10_6_0_V(reg_bend[10][6][0]),
.bend_10_6_1_V(reg_bend[10][6][1]),
.bend_10_7_0_V(reg_bend[10][7][0]),
.bend_10_7_1_V(reg_bend[10][7][1]),
.bend_10_8_0_V(reg_bend[10][8][0]),
.bend_10_8_1_V(reg_bend[10][8][1]),
.bend_11_0_0_V(reg_bend[11][0][0]),
.bend_11_0_1_V(reg_bend[11][0][1]),
.bend_11_1_0_V(reg_bend[11][1][0]),
.bend_11_1_1_V(reg_bend[11][1][1]),
.bend_11_2_0_V(reg_bend[11][2][0]),
.bend_11_2_1_V(reg_bend[11][2][1]),
.bend_11_3_0_V(reg_bend[11][3][0]),
.bend_11_3_1_V(reg_bend[11][3][1]),
.bend_11_4_0_V(reg_bend[11][4][0]),
.bend_11_4_1_V(reg_bend[11][4][1]),
.bend_11_5_0_V(reg_bend[11][5][0]),
.bend_11_5_1_V(reg_bend[11][5][1]),
.bend_11_6_0_V(reg_bend[11][6][0]),
.bend_11_6_1_V(reg_bend[11][6][1]),
.bend_11_7_0_V(reg_bend[11][7][0]),
.bend_11_7_1_V(reg_bend[11][7][1]),
.bend_11_8_0_V(reg_bend[11][8][0]),
.bend_11_8_1_V(reg_bend[11][8][1]),
.cs_0_V(reg_cs[0]),
.cs_1_V(reg_cs[1]),
.cs_2_V(reg_cs[2]),
.cs_3_V(reg_cs[3]),
.cs_4_V(reg_cs[4]),
.cs_5_V(reg_cs[5]),
.endcap_V(reg_endcap),
.sector_V(reg_sector),
.lat_test_V(reg_lat_test),
.core_config_V(reg_core_config),
.r_in_V(reg_r_in),
.we_V(reg_we),
.addr_V(reg_addr),
.sel_V(reg_sel),
.model_out_0_V(wire_model_out[0]),
.model_out_1_V(wire_model_out[1]),
.model_out_2_V(wire_model_out[2]),
.model_out_3_V(wire_model_out[3]),
.model_out_4_V(wire_model_out[4]),
.model_out_5_V(wire_model_out[5]),
.model_out_6_V(wire_model_out[6]),
.model_out_7_V(wire_model_out[7]),
.model_out_8_V(wire_model_out[8]),
.model_out_9_V(wire_model_out[9]),
.model_out_10_V(wire_model_out[10]),
.model_out_11_V(wire_model_out[11]),
.model_out_12_V(wire_model_out[12]),
.model_out_13_V(wire_model_out[13]),
.model_out_14_V(wire_model_out[14]),
.model_out_15_V(wire_model_out[15]),
.model_out_16_V(wire_model_out[16]),
.model_out_17_V(wire_model_out[17]),
.model_out_18_V(wire_model_out[18]),
.model_out_19_V(wire_model_out[19]),
.model_out_20_V(wire_model_out[20]),
.model_out_21_V(wire_model_out[21]),
.model_out_22_V(wire_model_out[22]),
.model_out_23_V(wire_model_out[23]),
.model_out_24_V(wire_model_out[24]),
.model_out_25_V(wire_model_out[25]),
.model_out_26_V(wire_model_out[26]),
.model_out_27_V(wire_model_out[27]),
.model_out_28_V(wire_model_out[28]),
.model_out_29_V(wire_model_out[29]),
.model_out_30_V(wire_model_out[30]),
.model_out_31_V(wire_model_out[31]),
.model_out_32_V(wire_model_out[32]),
.model_out_33_V(wire_model_out[33]),
.model_out_34_V(wire_model_out[34]),
.model_out_35_V(wire_model_out[35]),
.model_out_36_V(wire_model_out[36]),
.model_out_37_V(wire_model_out[37]),
.model_out_38_V(wire_model_out[38]),
.model_out_39_V(wire_model_out[39]),
.model_out_40_V(wire_model_out[40]),
.model_out_41_V(wire_model_out[41]),
.model_out_42_V(wire_model_out[42]),
.model_out_43_V(wire_model_out[43]),
.model_out_44_V(wire_model_out[44]),
.model_out_45_V(wire_model_out[45]),
.model_out_46_V(wire_model_out[46]),
.model_out_47_V(wire_model_out[47]),
.model_out_48_V(wire_model_out[48]),
.model_out_49_V(wire_model_out[49]),
.model_out_50_V(wire_model_out[50]),
.model_out_51_V(wire_model_out[51]),
.model_out_52_V(wire_model_out[52]),
.model_out_53_V(wire_model_out[53]),
.model_out_54_V(wire_model_out[54]),
.model_out_55_V(wire_model_out[55]),
.model_out_56_V(wire_model_out[56]),
.model_out_57_V(wire_model_out[57]),
.model_out_58_V(wire_model_out[58]),
.model_out_59_V(wire_model_out[59]),
.model_out_60_V(wire_model_out[60]),
.model_out_61_V(wire_model_out[61]),
.model_out_62_V(wire_model_out[62]),
.model_out_63_V(wire_model_out[63]),
.model_out_64_V(wire_model_out[64]),
.model_out_65_V(wire_model_out[65]),
.model_out_66_V(wire_model_out[66]),
.model_out_67_V(wire_model_out[67]),
.model_out_68_V(wire_model_out[68]),
.model_out_69_V(wire_model_out[69]),
.model_out_70_V(wire_model_out[70]),
.model_out_71_V(wire_model_out[71]),
.model_out_72_V(wire_model_out[72]),
.model_out_73_V(wire_model_out[73]),
.model_out_74_V(wire_model_out[74]),
.model_out_75_V(wire_model_out[75]),
.model_out_76_V(wire_model_out[76]),
.model_out_77_V(wire_model_out[77]),
.model_out_78_V(wire_model_out[78]),
.model_out_79_V(wire_model_out[79]),
.model_out_80_V(wire_model_out[80]),
.model_out_81_V(wire_model_out[81]),
.model_out_82_V(wire_model_out[82]),
.model_out_83_V(wire_model_out[83]),
.model_out_84_V(wire_model_out[84]),
.model_out_85_V(wire_model_out[85]),
.model_out_86_V(wire_model_out[86]),
.model_out_87_V(wire_model_out[87]),
.model_out_88_V(wire_model_out[88]),
.model_out_89_V(wire_model_out[89]),
.model_out_90_V(wire_model_out[90]),
.model_out_91_V(wire_model_out[91]),
.model_out_92_V(wire_model_out[92]),
.model_out_93_V(wire_model_out[93]),
.model_out_94_V(wire_model_out[94]),
.model_out_95_V(wire_model_out[95]),
.model_out_96_V(wire_model_out[96]),
.model_out_97_V(wire_model_out[97]),
.model_out_98_V(wire_model_out[98]),
.model_out_99_V(wire_model_out[99]),
.model_out_100_V(wire_model_out[100]),
.model_out_101_V(wire_model_out[101]),
.model_out_102_V(wire_model_out[102]),
.model_out_103_V(wire_model_out[103]),
.model_out_104_V(wire_model_out[104]),
.model_out_105_V(wire_model_out[105]),
.model_out_106_V(wire_model_out[106]),
.model_out_107_V(wire_model_out[107]),
.model_out_108_V(wire_model_out[108]),
.model_out_109_V(wire_model_out[109]),
.model_out_110_V(wire_model_out[110]),
.model_out_111_V(wire_model_out[111]),
.model_out_112_V(wire_model_out[112]),
.model_out_113_V(wire_model_out[113]),
.model_out_114_V(wire_model_out[114]),
.model_out_115_V(wire_model_out[115]),
.model_out_116_V(wire_model_out[116]),
.model_out_117_V(wire_model_out[117]),
.model_out_118_V(wire_model_out[118]),
.model_out_119_V(wire_model_out[119]),
.model_out_120_V(wire_model_out[120]),
.model_out_121_V(wire_model_out[121]),
.model_out_122_V(wire_model_out[122]),
.model_out_123_V(wire_model_out[123]),
.model_out_124_V(wire_model_out[124]),
.model_out_125_V(wire_model_out[125]),
.model_out_126_V(wire_model_out[126]),
.model_out_127_V(wire_model_out[127]),
.model_out_128_V(wire_model_out[128]),
.model_out_129_V(wire_model_out[129]),
.model_out_130_V(wire_model_out[130]),
.model_out_131_V(wire_model_out[131]),
.model_out_132_V(wire_model_out[132]),
.model_out_133_V(wire_model_out[133]),
.model_out_134_V(wire_model_out[134]),
.model_out_135_V(wire_model_out[135]),
.model_out_136_V(wire_model_out[136]),
.model_out_137_V(wire_model_out[137]),
.model_out_138_V(wire_model_out[138]),
.model_out_139_V(wire_model_out[139]),
.model_out_140_V(wire_model_out[140]),
.model_out_141_V(wire_model_out[141]),
.model_out_142_V(wire_model_out[142]),
.model_out_143_V(wire_model_out[143]),
.model_out_144_V(wire_model_out[144]),
.model_out_145_V(wire_model_out[145]),
.model_out_146_V(wire_model_out[146]),
.model_out_147_V(wire_model_out[147]),
.model_out_148_V(wire_model_out[148]),
.model_out_149_V(wire_model_out[149]),
.model_out_150_V(wire_model_out[150]),
.model_out_151_V(wire_model_out[151]),
.model_out_152_V(wire_model_out[152]),
.model_out_153_V(wire_model_out[153]),
.model_out_154_V(wire_model_out[154]),
.model_out_155_V(wire_model_out[155]),
.model_out_156_V(wire_model_out[156]),
.model_out_157_V(wire_model_out[157]),
.model_out_158_V(wire_model_out[158]),
.model_out_159_V(wire_model_out[159]),
.model_out_160_V(wire_model_out[160]),
.model_out_161_V(wire_model_out[161]),
.model_out_162_V(wire_model_out[162]),
.model_out_163_V(wire_model_out[163]),
.model_out_164_V(wire_model_out[164]),
.model_out_165_V(wire_model_out[165]),
.model_out_166_V(wire_model_out[166]),
.model_out_167_V(wire_model_out[167]),
.model_out_168_V(wire_model_out[168]),
.model_out_169_V(wire_model_out[169]),
.model_out_170_V(wire_model_out[170]),
.model_out_171_V(wire_model_out[171]),
.model_out_172_V(wire_model_out[172]),
.model_out_173_V(wire_model_out[173]),
.model_out_174_V(wire_model_out[174]),
.model_out_175_V(wire_model_out[175]),
.model_out_176_V(wire_model_out[176]),
.model_out_177_V(wire_model_out[177]),
.model_out_178_V(wire_model_out[178]),
.model_out_179_V(wire_model_out[179]),
.model_out_180_V(wire_model_out[180]),
.model_out_181_V(wire_model_out[181]),
.model_out_182_V(wire_model_out[182]),
.model_out_183_V(wire_model_out[183]),
.model_out_184_V(wire_model_out[184]),
.model_out_185_V(wire_model_out[185]),
.model_out_186_V(wire_model_out[186]),
.model_out_187_V(wire_model_out[187]),
.model_out_188_V(wire_model_out[188]),
.model_out_189_V(wire_model_out[189]),
.model_out_190_V(wire_model_out[190]),
.model_out_191_V(wire_model_out[191]),
.model_out_192_V(wire_model_out[192]),
.model_out_193_V(wire_model_out[193]),
.model_out_194_V(wire_model_out[194]),
.model_out_195_V(wire_model_out[195]),
.model_out_196_V(wire_model_out[196]),
.model_out_197_V(wire_model_out[197]),
.model_out_198_V(wire_model_out[198]),
.model_out_199_V(wire_model_out[199]),
.model_out_200_V(wire_model_out[200]),
.model_out_201_V(wire_model_out[201]),
.model_out_202_V(wire_model_out[202]),
.model_out_203_V(wire_model_out[203]),
.model_out_204_V(wire_model_out[204]),
.model_out_205_V(wire_model_out[205]),
.model_out_206_V(wire_model_out[206]),
.model_out_207_V(wire_model_out[207]),
.model_out_208_V(wire_model_out[208]),
.model_out_209_V(wire_model_out[209]),
.model_out_210_V(wire_model_out[210]),
.model_out_211_V(wire_model_out[211]),
.model_out_212_V(wire_model_out[212]),
.model_out_213_V(wire_model_out[213]),
.model_out_214_V(wire_model_out[214]),
.model_out_215_V(wire_model_out[215]),
.r_out_V(wire_r_out),
.model_out_0_V_ap_vld(),
.model_out_1_V_ap_vld(),
.model_out_2_V_ap_vld(),
.model_out_3_V_ap_vld(),
.model_out_4_V_ap_vld(),
.model_out_5_V_ap_vld(),
.model_out_6_V_ap_vld(),
.model_out_7_V_ap_vld(),
.model_out_8_V_ap_vld(),
.model_out_9_V_ap_vld(),
.model_out_10_V_ap_vld(),
.model_out_11_V_ap_vld(),
.model_out_12_V_ap_vld(),
.model_out_13_V_ap_vld(),
.model_out_14_V_ap_vld(),
.model_out_15_V_ap_vld(),
.model_out_16_V_ap_vld(),
.model_out_17_V_ap_vld(),
.model_out_18_V_ap_vld(),
.model_out_19_V_ap_vld(),
.model_out_20_V_ap_vld(),
.model_out_21_V_ap_vld(),
.model_out_22_V_ap_vld(),
.model_out_23_V_ap_vld(),
.model_out_24_V_ap_vld(),
.model_out_25_V_ap_vld(),
.model_out_26_V_ap_vld(),
.model_out_27_V_ap_vld(),
.model_out_28_V_ap_vld(),
.model_out_29_V_ap_vld(),
.model_out_30_V_ap_vld(),
.model_out_31_V_ap_vld(),
.model_out_32_V_ap_vld(),
.model_out_33_V_ap_vld(),
.model_out_34_V_ap_vld(),
.model_out_35_V_ap_vld(),
.model_out_36_V_ap_vld(),
.model_out_37_V_ap_vld(),
.model_out_38_V_ap_vld(),
.model_out_39_V_ap_vld(),
.model_out_40_V_ap_vld(),
.model_out_41_V_ap_vld(),
.model_out_42_V_ap_vld(),
.model_out_43_V_ap_vld(),
.model_out_44_V_ap_vld(),
.model_out_45_V_ap_vld(),
.model_out_46_V_ap_vld(),
.model_out_47_V_ap_vld(),
.model_out_48_V_ap_vld(),
.model_out_49_V_ap_vld(),
.model_out_50_V_ap_vld(),
.model_out_51_V_ap_vld(),
.model_out_52_V_ap_vld(),
.model_out_53_V_ap_vld(),
.model_out_54_V_ap_vld(),
.model_out_55_V_ap_vld(),
.model_out_56_V_ap_vld(),
.model_out_57_V_ap_vld(),
.model_out_58_V_ap_vld(),
.model_out_59_V_ap_vld(),
.model_out_60_V_ap_vld(),
.model_out_61_V_ap_vld(),
.model_out_62_V_ap_vld(),
.model_out_63_V_ap_vld(),
.model_out_64_V_ap_vld(),
.model_out_65_V_ap_vld(),
.model_out_66_V_ap_vld(),
.model_out_67_V_ap_vld(),
.model_out_68_V_ap_vld(),
.model_out_69_V_ap_vld(),
.model_out_70_V_ap_vld(),
.model_out_71_V_ap_vld(),
.model_out_72_V_ap_vld(),
.model_out_73_V_ap_vld(),
.model_out_74_V_ap_vld(),
.model_out_75_V_ap_vld(),
.model_out_76_V_ap_vld(),
.model_out_77_V_ap_vld(),
.model_out_78_V_ap_vld(),
.model_out_79_V_ap_vld(),
.model_out_80_V_ap_vld(),
.model_out_81_V_ap_vld(),
.model_out_82_V_ap_vld(),
.model_out_83_V_ap_vld(),
.model_out_84_V_ap_vld(),
.model_out_85_V_ap_vld(),
.model_out_86_V_ap_vld(),
.model_out_87_V_ap_vld(),
.model_out_88_V_ap_vld(),
.model_out_89_V_ap_vld(),
.model_out_90_V_ap_vld(),
.model_out_91_V_ap_vld(),
.model_out_92_V_ap_vld(),
.model_out_93_V_ap_vld(),
.model_out_94_V_ap_vld(),
.model_out_95_V_ap_vld(),
.model_out_96_V_ap_vld(),
.model_out_97_V_ap_vld(),
.model_out_98_V_ap_vld(),
.model_out_99_V_ap_vld(),
.model_out_100_V_ap_vld(),
.model_out_101_V_ap_vld(),
.model_out_102_V_ap_vld(),
.model_out_103_V_ap_vld(),
.model_out_104_V_ap_vld(),
.model_out_105_V_ap_vld(),
.model_out_106_V_ap_vld(),
.model_out_107_V_ap_vld(),
.model_out_108_V_ap_vld(),
.model_out_109_V_ap_vld(),
.model_out_110_V_ap_vld(),
.model_out_111_V_ap_vld(),
.model_out_112_V_ap_vld(),
.model_out_113_V_ap_vld(),
.model_out_114_V_ap_vld(),
.model_out_115_V_ap_vld(),
.model_out_116_V_ap_vld(),
.model_out_117_V_ap_vld(),
.model_out_118_V_ap_vld(),
.model_out_119_V_ap_vld(),
.model_out_120_V_ap_vld(),
.model_out_121_V_ap_vld(),
.model_out_122_V_ap_vld(),
.model_out_123_V_ap_vld(),
.model_out_124_V_ap_vld(),
.model_out_125_V_ap_vld(),
.model_out_126_V_ap_vld(),
.model_out_127_V_ap_vld(),
.model_out_128_V_ap_vld(),
.model_out_129_V_ap_vld(),
.model_out_130_V_ap_vld(),
.model_out_131_V_ap_vld(),
.model_out_132_V_ap_vld(),
.model_out_133_V_ap_vld(),
.model_out_134_V_ap_vld(),
.model_out_135_V_ap_vld(),
.model_out_136_V_ap_vld(),
.model_out_137_V_ap_vld(),
.model_out_138_V_ap_vld(),
.model_out_139_V_ap_vld(),
.model_out_140_V_ap_vld(),
.model_out_141_V_ap_vld(),
.model_out_142_V_ap_vld(),
.model_out_143_V_ap_vld(),
.model_out_144_V_ap_vld(),
.model_out_145_V_ap_vld(),
.model_out_146_V_ap_vld(),
.model_out_147_V_ap_vld(),
.model_out_148_V_ap_vld(),
.model_out_149_V_ap_vld(),
.model_out_150_V_ap_vld(),
.model_out_151_V_ap_vld(),
.model_out_152_V_ap_vld(),
.model_out_153_V_ap_vld(),
.model_out_154_V_ap_vld(),
.model_out_155_V_ap_vld(),
.model_out_156_V_ap_vld(),
.model_out_157_V_ap_vld(),
.model_out_158_V_ap_vld(),
.model_out_159_V_ap_vld(),
.model_out_160_V_ap_vld(),
.model_out_161_V_ap_vld(),
.model_out_162_V_ap_vld(),
.model_out_163_V_ap_vld(),
.model_out_164_V_ap_vld(),
.model_out_165_V_ap_vld(),
.model_out_166_V_ap_vld(),
.model_out_167_V_ap_vld(),
.model_out_168_V_ap_vld(),
.model_out_169_V_ap_vld(),
.model_out_170_V_ap_vld(),
.model_out_171_V_ap_vld(),
.model_out_172_V_ap_vld(),
.model_out_173_V_ap_vld(),
.model_out_174_V_ap_vld(),
.model_out_175_V_ap_vld(),
.model_out_176_V_ap_vld(),
.model_out_177_V_ap_vld(),
.model_out_178_V_ap_vld(),
.model_out_179_V_ap_vld(),
.model_out_180_V_ap_vld(),
.model_out_181_V_ap_vld(),
.model_out_182_V_ap_vld(),
.model_out_183_V_ap_vld(),
.model_out_184_V_ap_vld(),
.model_out_185_V_ap_vld(),
.model_out_186_V_ap_vld(),
.model_out_187_V_ap_vld(),
.model_out_188_V_ap_vld(),
.model_out_189_V_ap_vld(),
.model_out_190_V_ap_vld(),
.model_out_191_V_ap_vld(),
.model_out_192_V_ap_vld(),
.model_out_193_V_ap_vld(),
.model_out_194_V_ap_vld(),
.model_out_195_V_ap_vld(),
.model_out_196_V_ap_vld(),
.model_out_197_V_ap_vld(),
.model_out_198_V_ap_vld(),
.model_out_199_V_ap_vld(),
.model_out_200_V_ap_vld(),
.model_out_201_V_ap_vld(),
.model_out_202_V_ap_vld(),
.model_out_203_V_ap_vld(),
.model_out_204_V_ap_vld(),
.model_out_205_V_ap_vld(),
.model_out_206_V_ap_vld(),
.model_out_207_V_ap_vld(),
.model_out_208_V_ap_vld(),
.model_out_209_V_ap_vld(),
.model_out_210_V_ap_vld(),
.model_out_211_V_ap_vld(),
.model_out_212_V_ap_vld(),
.model_out_213_V_ap_vld(),
.model_out_214_V_ap_vld(),
.model_out_215_V_ap_vld()
    );

    integer i;
    integer j;
    integer k;
    integer l;

    always @(posedge clock) begin
        if (reset == 1'h1) begin

// RESET LOGIC

for (i=0; i<12; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		reg_vpf[i][j] <= 0;
	end
end
for (i=0; i<12; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_q[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_wg[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_hstr[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_cpat[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_ph_rpc[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_th_rpc[i][j][k] <= 0;
		end
	end
end
for (i=0; i<12; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_time[i][j][k] <= 0;
		end
	end
end
for (i=0; i<12; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_bend[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	reg_cs[i] <= 0;
end
reg_endcap <= 0;
reg_sector <= 0;
reg_lat_test <= 0;
reg_core_config <= 0;
reg_r_in <= 0;
reg_we <= 0;
reg_addr <= 0;
reg_sel <= 0;
for (i=0; i<216; i=i+1) begin
	reg_model_out[i] <= 0;
end
bus_model_out <= 0;
reg_r_out <= 0;
bus_r_out <= 0;
        end else begin

// SHIFT LOGIC


// SHIFT LOGIC - INPUT: [vpf]

if (feed_in_vpf == 1'h1) begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			if (j==0) begin
				if (i==0) begin
					reg_vpf[i][j] <= bus_vpf;
				end else begin
					reg_vpf[i][j] <= reg_vpf[i-1][9-1];
				end
			end else begin
				reg_vpf[i][j] <= reg_vpf[i][j-1];
			end
		end
	end
end else begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			reg_vpf[i][j] <= reg_vpf[i][j];
		end
	end
end

// SHIFT LOGIC - INPUT: [q]

if (feed_in_q == 1'h1) begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_q[i][j][k] <= bus_q;
						end else begin
							reg_q[i][j][k] <= reg_q[i-1][9-1][2-1];
						end
					end else begin
						reg_q[i][j][k] <= reg_q[i][j-1][2-1];
					end
				end else begin
					reg_q[i][j][k] <= reg_q[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_q[i][j][k] <= reg_q[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [wg]

if (feed_in_wg == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_wg[i][j][k] <= bus_wg;
						end else begin
							reg_wg[i][j][k] <= reg_wg[i-1][9-1][2-1];
						end
					end else begin
						reg_wg[i][j][k] <= reg_wg[i][j-1][2-1];
					end
				end else begin
					reg_wg[i][j][k] <= reg_wg[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_wg[i][j][k] <= reg_wg[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [hstr]

if (feed_in_hstr == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_hstr[i][j][k] <= bus_hstr;
						end else begin
							reg_hstr[i][j][k] <= reg_hstr[i-1][9-1][2-1];
						end
					end else begin
						reg_hstr[i][j][k] <= reg_hstr[i][j-1][2-1];
					end
				end else begin
					reg_hstr[i][j][k] <= reg_hstr[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_hstr[i][j][k] <= reg_hstr[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [cpat]

if (feed_in_cpat == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_cpat[i][j][k] <= bus_cpat;
						end else begin
							reg_cpat[i][j][k] <= reg_cpat[i-1][9-1][2-1];
						end
					end else begin
						reg_cpat[i][j][k] <= reg_cpat[i][j-1][2-1];
					end
				end else begin
					reg_cpat[i][j][k] <= reg_cpat[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_cpat[i][j][k] <= reg_cpat[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [ph_rpc]

if (feed_in_ph_rpc == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_ph_rpc[i][j][k] <= bus_ph_rpc;
						end else begin
							reg_ph_rpc[i][j][k] <= reg_ph_rpc[i-1][9-1][2-1];
						end
					end else begin
						reg_ph_rpc[i][j][k] <= reg_ph_rpc[i][j-1][2-1];
					end
				end else begin
					reg_ph_rpc[i][j][k] <= reg_ph_rpc[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_ph_rpc[i][j][k] <= reg_ph_rpc[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [th_rpc]

if (feed_in_th_rpc == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_th_rpc[i][j][k] <= bus_th_rpc;
						end else begin
							reg_th_rpc[i][j][k] <= reg_th_rpc[i-1][9-1][2-1];
						end
					end else begin
						reg_th_rpc[i][j][k] <= reg_th_rpc[i][j-1][2-1];
					end
				end else begin
					reg_th_rpc[i][j][k] <= reg_th_rpc[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_th_rpc[i][j][k] <= reg_th_rpc[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [time]

if (feed_in_time == 1'h1) begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_time[i][j][k] <= bus_time;
						end else begin
							reg_time[i][j][k] <= reg_time[i-1][9-1][2-1];
						end
					end else begin
						reg_time[i][j][k] <= reg_time[i][j-1][2-1];
					end
				end else begin
					reg_time[i][j][k] <= reg_time[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_time[i][j][k] <= reg_time[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [bend]

if (feed_in_bend == 1'h1) begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_bend[i][j][k] <= bus_bend;
						end else begin
							reg_bend[i][j][k] <= reg_bend[i-1][9-1][2-1];
						end
					end else begin
						reg_bend[i][j][k] <= reg_bend[i][j-1][2-1];
					end
				end else begin
					reg_bend[i][j][k] <= reg_bend[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<12; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_bend[i][j][k] <= reg_bend[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [cs]

if (feed_in_cs == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		if (i==0) begin
			reg_cs[i] <= bus_cs;
		end else begin
			reg_cs[i] <= reg_cs[i-1];
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		reg_cs[i] <= reg_cs[i];
	end
end

// SHIFT LOGIC - INPUT: [endcap]

if (feed_in_endcap == 1'h1) begin
	reg_endcap <= bus_endcap;
end else begin
	reg_endcap <= reg_endcap;
end

// SHIFT LOGIC - INPUT: [sector]

if (feed_in_sector == 1'h1) begin
	reg_sector <= bus_sector;
end else begin
	reg_sector <= reg_sector;
end

// SHIFT LOGIC - INPUT: [lat_test]

if (feed_in_lat_test == 1'h1) begin
	reg_lat_test <= bus_lat_test;
end else begin
	reg_lat_test <= reg_lat_test;
end

// SHIFT LOGIC - INPUT: [core_config]

if (feed_in_core_config == 1'h1) begin
	reg_core_config <= bus_core_config;
end else begin
	reg_core_config <= reg_core_config;
end

// SHIFT LOGIC - INPUT: [r_in]

if (feed_in_r_in == 1'h1) begin
	reg_r_in <= bus_r_in;
end else begin
	reg_r_in <= reg_r_in;
end

// SHIFT LOGIC - INPUT: [we]

if (feed_in_we == 1'h1) begin
	reg_we <= bus_we;
end else begin
	reg_we <= reg_we;
end

// SHIFT LOGIC - INPUT: [addr]

if (feed_in_addr == 1'h1) begin
	reg_addr <= bus_addr;
end else begin
	reg_addr <= reg_addr;
end

// SHIFT LOGIC - INPUT: [sel]

if (feed_in_sel == 1'h1) begin
	reg_sel <= bus_sel;
end else begin
	reg_sel <= reg_sel;
end

// SHIFT LOGIC - OUTPUT: [model_out]

if (feed_out_model_out == 1'h1) begin
	for (i=0; i<216; i=i+1) begin
		if (i==0) begin
			reg_model_out[i] <= bus_model_out;
		end else begin
			reg_model_out[i] <= reg_model_out[i-1];
			if (i==216-1) begin
				bus_model_out <= reg_model_out[i];
			end
		end
	end
end else if (load_out_model_out == 1'h1) begin
	for (i=0; i<216; i=i+1) begin
		reg_model_out[i] <= wire_model_out[i];
	end
end else begin
	for (i=0; i<216; i=i+1) begin
		reg_model_out[i] <= reg_model_out[i];
	end
	bus_model_out <= bus_model_out;
end

// SHIFT LOGIC - OUTPUT: [r_out]

if (feed_out_r_out == 1'h1) begin
	bus_r_out <= reg_r_out;
end else if (load_out_r_out == 1'h1) begin
	reg_r_out <= wire_r_out;
end else begin
	reg_r_out <= reg_r_out;
	bus_r_out <= bus_r_out;
end
        end
    end

endmodule
